/* This file is just an example for PRVTDNN, use Chisel to generate your
* version*/
module LoadWeightBias(
  input         clock,
  input         reset,
  input  [15:0] io_bramIF_wrData,
  output [15:0] io_bramIF_rdData,
  input  [8:0]  io_bramIF_wrAddr,
  input  [8:0]  io_bramIF_rdAddr,
  input         io_bramIF_wrEn,
  output [15:0] io_outWeight_0,
  output [15:0] io_outWeight_1,
  output [15:0] io_outWeight_2,
  output [15:0] io_outWeight_3,
  output [15:0] io_outWeight_4,
  output [15:0] io_outWeight_5,
  output [15:0] io_outWeight_6,
  output [15:0] io_outWeight_7,
  output [15:0] io_outWeight_8,
  output [15:0] io_outWeight_9,
  output [15:0] io_outBias_0,
  output [15:0] io_outBias_1,
  output [15:0] io_outBias_2,
  output [15:0] io_outBias_3,
  output [15:0] io_outBias_4,
  output [15:0] io_outBias_5,
  output [15:0] io_outBias_6,
  output [15:0] io_outBias_7,
  output [15:0] io_outBias_8,
  output [15:0] io_outBias_9,
  output [2:0]  io_outWtValid,
  output [2:0]  io_outBiasValid,
  input         io_load
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_GARBAGE_ASSIGN
  reg [15:0] mem [0:407]; // @[LoadWeightBias.scala 42:26]
  wire  mem_io_bramIF_rdData_MPORT_en; // @[LoadWeightBias.scala 42:26]
  wire [8:0] mem_io_bramIF_rdData_MPORT_addr; // @[LoadWeightBias.scala 42:26]
  wire [15:0] mem_io_bramIF_rdData_MPORT_data; // @[LoadWeightBias.scala 42:26]
  wire  mem_memRdDataWire_MPORT_en; // @[LoadWeightBias.scala 42:26]
  wire [8:0] mem_memRdDataWire_MPORT_addr; // @[LoadWeightBias.scala 42:26]
  wire [15:0] mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 42:26]
  wire  mem_memRdDataWire_MPORT_1_en; // @[LoadWeightBias.scala 42:26]
  wire [8:0] mem_memRdDataWire_MPORT_1_addr; // @[LoadWeightBias.scala 42:26]
  wire [15:0] mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 42:26]
  wire [15:0] mem_MPORT_data; // @[LoadWeightBias.scala 42:26]
  wire [8:0] mem_MPORT_addr; // @[LoadWeightBias.scala 42:26]
  wire  mem_MPORT_mask; // @[LoadWeightBias.scala 42:26]
  wire  mem_MPORT_en; // @[LoadWeightBias.scala 42:26]
  reg  mem_io_bramIF_rdData_MPORT_en_pipe_0;
  reg [8:0] mem_io_bramIF_rdData_MPORT_addr_pipe_0;
  reg  mem_memRdDataWire_MPORT_en_pipe_0;
  reg [8:0] mem_memRdDataWire_MPORT_addr_pipe_0;
  reg  mem_memRdDataWire_MPORT_1_en_pipe_0;
  reg [8:0] mem_memRdDataWire_MPORT_1_addr_pipe_0;
  reg [2:0] wtValidReg; // @[LoadWeightBias.scala 56:26]
  reg [2:0] biasValidReg; // @[LoadWeightBias.scala 57:26]
  reg [1:0] layerCnt_value; // @[Counter.scala 61:40]
  reg [4:0] rowCnt_value; // @[Counter.scala 61:40]
  reg [3:0] columnCnt_value; // @[Counter.scala 61:40]
  reg [15:0] weightReg_0; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_1; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_2; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_3; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_4; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_5; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_6; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_7; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_8; // @[LoadWeightBias.scala 62:26]
  reg [15:0] weightReg_9; // @[LoadWeightBias.scala 62:26]
  reg [15:0] biasReg_0; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_1; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_2; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_3; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_4; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_5; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_6; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_7; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_8; // @[LoadWeightBias.scala 63:26]
  reg [15:0] biasReg_9; // @[LoadWeightBias.scala 63:26]
  reg [1:0] stateReg; // @[LoadWeightBias.scala 68:30]
  reg [8:0] addrReg; // @[LoadWeightBias.scala 69:30]
  reg  loadWFinReg; // @[LoadWeightBias.scala 70:43]
  reg  loadBFinReg; // @[LoadWeightBias.scala 70:43]
  wire [1:0] _GEN_11 = loadBFinReg ? 2'h0 : 2'h2; // @[LoadWeightBias.scala 82:{33,44} 83:44]
  wire  _switchFlagW_T = layerCnt_value == 2'h2; // @[LoadWeightBias.scala 94:36]
  wire [4:0] _GEN_16 = 2'h1 == layerCnt_value ? 5'ha : 5'h14; // @[LoadWeightBias.scala 95:{56,56}]
  wire [4:0] _GEN_17 = 2'h2 == layerCnt_value ? 5'ha : _GEN_16; // @[LoadWeightBias.scala 95:{56,56}]
  wire [4:0] _switchFlagW_T_2 = _GEN_17 - 5'h1; // @[LoadWeightBias.scala 95:56]
  wire  _switchFlagW_T_3 = rowCnt_value == _switchFlagW_T_2; // @[LoadWeightBias.scala 95:27]
  wire  _switchFlagW_T_4 = layerCnt_value == 2'h2 & _switchFlagW_T_3; // @[LoadWeightBias.scala 94:56]
  wire [3:0] _GEN_20 = 2'h2 == layerCnt_value ? 4'h8 : 4'ha; // @[LoadWeightBias.scala 96:{62,62}]
  wire [3:0] _switchFlagW_T_6 = _GEN_20 - 4'h1; // @[LoadWeightBias.scala 96:62]
  wire  _switchFlagW_T_7 = columnCnt_value == _switchFlagW_T_6; // @[LoadWeightBias.scala 96:30]
  wire  switchFlagW = _switchFlagW_T_4 & _switchFlagW_T_7; // @[LoadWeightBias.scala 95:62]
  wire  switchFlagB = _switchFlagW_T & _switchFlagW_T_7; // @[LoadWeightBias.scala 98:56]
  wire  _T_3 = stateReg == 2'h0; // @[LoadWeightBias.scala 102:19]
  wire [8:0] _memRdDataWire_T_3 = addrReg + 9'h1; // @[LoadWeightBias.scala 106:43]
  wire  _T_5 = switchFlagW | loadWFinReg; // @[LoadWeightBias.scala 112:26]
  wire  _T_12 = _switchFlagW_T_3 & _switchFlagW_T_7; // @[LoadWeightBias.scala 119:67]
  wire [1:0] _value_T_1 = layerCnt_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _GEN_32 = _switchFlagW_T ? 2'h0 : _value_T_1; // @[Counter.scala 77:15 87:{20,28}]
  wire  wrap_1 = rowCnt_value == 5'h13; // @[Counter.scala 73:24]
  wire [4:0] _value_T_3 = rowCnt_value + 5'h1; // @[Counter.scala 77:24]
  wire [4:0] _GEN_33 = wrap_1 ? 5'h0 : _value_T_3; // @[Counter.scala 77:15 87:{20,28}]
  wire  wrap_2 = columnCnt_value == 4'h9; // @[Counter.scala 73:24]
  wire [3:0] _value_T_5 = columnCnt_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _GEN_34 = wrap_2 ? 4'h0 : _value_T_5; // @[Counter.scala 77:15 87:{20,28}]
  wire [4:0] _GEN_35 = _switchFlagW_T_7 ? _GEN_33 : rowCnt_value; // @[LoadWeightBias.scala 125:75 Counter.scala 61:40]
  wire [3:0] _GEN_36 = _switchFlagW_T_7 ? 4'h0 : _GEN_34; // @[LoadWeightBias.scala 125:75 Counter.scala 98:11]
  wire [3:0] _wtValidReg_T = 4'h1 << layerCnt_value; // @[OneHot.scala 57:35]
  wire [3:0] _GEN_65 = _switchFlagW_T_7 ? _wtValidReg_T : 4'h0; // @[LoadWeightBias.scala 137:67 138:24 140:24]
  wire [1:0] _GEN_68 = _switchFlagW_T_7 ? _GEN_32 : layerCnt_value; // @[LoadWeightBias.scala 148:71 Counter.scala 61:40]
  wire  _GEN_70 = switchFlagB | loadBFinReg; // @[LoadWeightBias.scala 144:26 145:25 70:43]
  wire  _GEN_85 = stateReg == 2'h2 & _GEN_70; // @[LoadWeightBias.scala 142:35 164:21]
  wire [3:0] _GEN_99 = stateReg == 2'h2 ? _GEN_65 : 4'h0; // @[LoadWeightBias.scala 142:35 171:22]
  wire  _GEN_100 = stateReg == 2'h2 & loadWFinReg; // @[LoadWeightBias.scala 142:35 163:21 70:43]
  wire [3:0] _GEN_112 = stateReg == 2'h1 ? 4'h0 : _GEN_99; // @[LoadWeightBias.scala 109:29 110:22]
  wire [3:0] _GEN_128 = stateReg == 2'h1 ? _GEN_65 : 4'h0; // @[LoadWeightBias.scala 109:29]
  assign mem_io_bramIF_rdData_MPORT_en = mem_io_bramIF_rdData_MPORT_en_pipe_0;
  assign mem_io_bramIF_rdData_MPORT_addr = mem_io_bramIF_rdData_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_io_bramIF_rdData_MPORT_data = mem[mem_io_bramIF_rdData_MPORT_addr]; // @[LoadWeightBias.scala 42:26]
  `else
  assign mem_io_bramIF_rdData_MPORT_data = mem_io_bramIF_rdData_MPORT_addr >= 9'h198 ? _RAND_0[15:0] :
    mem[mem_io_bramIF_rdData_MPORT_addr]; // @[LoadWeightBias.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_memRdDataWire_MPORT_en = mem_memRdDataWire_MPORT_en_pipe_0;
  assign mem_memRdDataWire_MPORT_addr = mem_memRdDataWire_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_memRdDataWire_MPORT_data = mem[mem_memRdDataWire_MPORT_addr]; // @[LoadWeightBias.scala 42:26]
  `else
  assign mem_memRdDataWire_MPORT_data = mem_memRdDataWire_MPORT_addr >= 9'h198 ? _RAND_1[15:0] :
    mem[mem_memRdDataWire_MPORT_addr]; // @[LoadWeightBias.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_memRdDataWire_MPORT_1_en = mem_memRdDataWire_MPORT_1_en_pipe_0;
  assign mem_memRdDataWire_MPORT_1_addr = mem_memRdDataWire_MPORT_1_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_memRdDataWire_MPORT_1_data = mem[mem_memRdDataWire_MPORT_1_addr]; // @[LoadWeightBias.scala 42:26]
  `else
  assign mem_memRdDataWire_MPORT_1_data = mem_memRdDataWire_MPORT_1_addr >= 9'h198 ? _RAND_2[15:0] :
    mem[mem_memRdDataWire_MPORT_1_addr]; // @[LoadWeightBias.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = io_bramIF_wrData;
  assign mem_MPORT_addr = io_bramIF_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_bramIF_wrEn;
  assign io_bramIF_rdData = mem_io_bramIF_rdData_MPORT_data; // @[LoadWeightBias.scala 48:22]
  assign io_outWeight_0 = weightReg_0; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_1 = weightReg_1; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_2 = weightReg_2; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_3 = weightReg_3; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_4 = weightReg_4; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_5 = weightReg_5; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_6 = weightReg_6; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_7 = weightReg_7; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_8 = weightReg_8; // @[LoadWeightBias.scala 175:21]
  assign io_outWeight_9 = weightReg_9; // @[LoadWeightBias.scala 175:21]
  assign io_outBias_0 = biasReg_0; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_1 = biasReg_1; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_2 = biasReg_2; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_3 = biasReg_3; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_4 = biasReg_4; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_5 = biasReg_5; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_6 = biasReg_6; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_7 = biasReg_7; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_8 = biasReg_8; // @[LoadWeightBias.scala 176:21]
  assign io_outBias_9 = biasReg_9; // @[LoadWeightBias.scala 176:21]
  assign io_outWtValid = wtValidReg; // @[LoadWeightBias.scala 177:21]
  assign io_outBiasValid = biasValidReg; // @[LoadWeightBias.scala 178:21]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[LoadWeightBias.scala 42:26]
    end
    mem_io_bramIF_rdData_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_bramIF_rdData_MPORT_addr_pipe_0 <= io_bramIF_rdAddr;
    end
    mem_memRdDataWire_MPORT_en_pipe_0 <= stateReg == 2'h0;
    if (stateReg == 2'h0) begin
      mem_memRdDataWire_MPORT_addr_pipe_0 <= 9'h0;
    end
    if (_T_3) begin
      mem_memRdDataWire_MPORT_1_en_pipe_0 <= 1'h0;
    end else begin
      mem_memRdDataWire_MPORT_1_en_pipe_0 <= 1'h1;
    end
    if (_T_3 ? 1'h0 : 1'h1) begin
      mem_memRdDataWire_MPORT_1_addr_pipe_0 <= addrReg + 9'h1;
    end
    wtValidReg <= _GEN_128[2:0];
    biasValidReg <= _GEN_112[2:0];
    if (reset) begin // @[Counter.scala 61:40]
      layerCnt_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (switchFlagW | loadWFinReg) begin // @[LoadWeightBias.scala 112:41]
        layerCnt_value <= 2'h0; // @[Counter.scala 98:11]
      end else if (_T_12) begin // @[LoadWeightBias.scala 120:75]
        layerCnt_value <= _GEN_32;
      end
    end else if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
      if (!(switchFlagB)) begin // @[LoadWeightBias.scala 144:26]
        layerCnt_value <= _GEN_68;
      end
    end else begin
      layerCnt_value <= 2'h0; // @[Counter.scala 98:11]
    end
    if (reset) begin // @[Counter.scala 61:40]
      rowCnt_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (switchFlagW | loadWFinReg) begin // @[LoadWeightBias.scala 112:41]
        rowCnt_value <= 5'h0; // @[Counter.scala 98:11]
      end else if (_T_12) begin // @[LoadWeightBias.scala 120:75]
        rowCnt_value <= 5'h0; // @[Counter.scala 98:11]
      end else begin
        rowCnt_value <= _GEN_35;
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      rowCnt_value <= 5'h0; // @[Counter.scala 98:11]
    end
    if (reset) begin // @[Counter.scala 61:40]
      columnCnt_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (switchFlagW | loadWFinReg) begin // @[LoadWeightBias.scala 112:41]
        columnCnt_value <= 4'h0; // @[Counter.scala 98:11]
      end else if (_T_12) begin // @[LoadWeightBias.scala 120:75]
        columnCnt_value <= 4'h0; // @[Counter.scala 98:11]
      end else begin
        columnCnt_value <= _GEN_36;
      end
    end else if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
      if (switchFlagB) begin // @[LoadWeightBias.scala 144:26]
        columnCnt_value <= 4'h0; // @[Counter.scala 98:11]
      end else begin
        columnCnt_value <= _GEN_36;
      end
    end else begin
      columnCnt_value <= 4'h0; // @[Counter.scala 98:11]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h0 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_0 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_0 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_0 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h1 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_1 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_1 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_1 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h2 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_2 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_2 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_2 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h3 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_3 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_3 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_3 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h4 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_4 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_4 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_4 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h5 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_5 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_5 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_5 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h6 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_6 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_6 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_6 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h7 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_7 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_7 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_7 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h8 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_8 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_8 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_8 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~loadWFinReg) begin // @[LoadWeightBias.scala 136:28]
        if (4'h9 == columnCnt_value) begin // @[LoadWeightBias.scala 136:56]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            weightReg_9 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            weightReg_9 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end
    end else if (!(stateReg == 2'h2)) begin // @[LoadWeightBias.scala 142:35]
      weightReg_9 <= 16'sh0; // @[LoadWeightBias.scala 165:25]
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h0 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_0 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_0 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_0 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h1 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_1 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_1 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_1 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h2 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_2 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_2 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_2 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h3 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_3 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_3 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_3 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h4 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_4 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_4 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_4 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h5 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_5 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_5 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_5 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h6 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_6 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_6 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_6 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h7 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_7 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_7 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_7 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h8 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_8 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_8 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_8 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
        if (4'h9 == columnCnt_value) begin // @[LoadWeightBias.scala 156:34]
          if (stateReg == 2'h0) begin // @[LoadWeightBias.scala 102:28]
            biasReg_9 <= mem_memRdDataWire_MPORT_data; // @[LoadWeightBias.scala 103:23]
          end else begin
            biasReg_9 <= mem_memRdDataWire_MPORT_1_data; // @[LoadWeightBias.scala 106:23]
          end
        end
      end else begin
        biasReg_9 <= 16'sh0; // @[LoadWeightBias.scala 166:23]
      end
    end
    if (reset) begin // @[LoadWeightBias.scala 68:30]
      stateReg <= 2'h0; // @[LoadWeightBias.scala 68:30]
    end else if (2'h0 == stateReg) begin // @[LoadWeightBias.scala 72:21]
      if (io_load) begin // @[LoadWeightBias.scala 74:33]
        stateReg <= 2'h1; // @[LoadWeightBias.scala 74:44]
      end else begin
        stateReg <= 2'h0; // @[LoadWeightBias.scala 75:44]
      end
    end else if (2'h1 == stateReg) begin // @[LoadWeightBias.scala 72:21]
      if (loadWFinReg) begin // @[LoadWeightBias.scala 78:33]
        stateReg <= 2'h2; // @[LoadWeightBias.scala 78:44]
      end else begin
        stateReg <= 2'h1; // @[LoadWeightBias.scala 79:44]
      end
    end else if (2'h2 == stateReg) begin // @[LoadWeightBias.scala 72:21]
      stateReg <= _GEN_11;
    end
    if (reset) begin // @[LoadWeightBias.scala 69:30]
      addrReg <= 9'h0; // @[LoadWeightBias.scala 69:30]
    end else if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      if (~switchFlagW) begin // @[LoadWeightBias.scala 134:28]
        addrReg <= _memRdDataWire_T_3; // @[LoadWeightBias.scala 134:38]
      end
    end else if (stateReg == 2'h2) begin // @[LoadWeightBias.scala 142:35]
      addrReg <= _memRdDataWire_T_3; // @[LoadWeightBias.scala 155:17]
    end else begin
      addrReg <= 9'h0; // @[LoadWeightBias.scala 172:17]
    end
    if (reset) begin // @[LoadWeightBias.scala 70:43]
      loadWFinReg <= 1'h0; // @[LoadWeightBias.scala 70:43]
    end else if (stateReg == 2'h1) begin // @[LoadWeightBias.scala 109:29]
      loadWFinReg <= _T_5;
    end else begin
      loadWFinReg <= _GEN_100;
    end
    if (reset) begin // @[LoadWeightBias.scala 70:43]
      loadBFinReg <= 1'h0; // @[LoadWeightBias.scala 70:43]
    end else if (!(stateReg == 2'h1)) begin // @[LoadWeightBias.scala 109:29]
      loadBFinReg <= _GEN_85;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_0 = {1{`RANDOM}};
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE(
  input         clock,
  input  [15:0] io_inAct,
  input  [39:0] io_inWtPS,
  output [39:0] io_outWtPS,
  output [15:0] io_outAct,
  input         io_inwtValid
);
  reg [15:0] weightReg; // @[PE.scala 20:26]
  reg [15:0] actReg; // @[PE.scala 21:26]
  reg [39:0] parSumReg; // @[PE.scala 22:26]
  wire [31:0] _parSumReg_T = $signed(weightReg) * $signed(actReg); // @[PE.scala 26:40]
  wire [39:0] _GEN_2 = {{8{_parSumReg_T[31]}},_parSumReg_T}; // @[PE.scala 26:28]
  wire [39:0] _GEN_0 = io_inwtValid ? $signed(io_inWtPS) : $signed({{24{weightReg[15]}},weightReg}); // @[PE.scala 30:31 31:21 34:21]
  assign io_outWtPS = io_inwtValid ? $signed({{24{weightReg[15]}},weightReg}) : $signed(parSumReg); // @[PE.scala 30:31 32:21 35:21]
  assign io_outAct = actReg; // @[PE.scala 27:15]
  always @(posedge clock) begin
    weightReg <= _GEN_0[15:0];
    actReg <= io_inAct; // @[PE.scala 24:15]
    parSumReg <= $signed(io_inWtPS) + $signed(_GEN_2); // @[PE.scala 26:28]
  end
endmodule
module SystolicArray(
  input         clock,
  input  [15:0] io_inAct_0,
  input  [15:0] io_inAct_1,
  input  [15:0] io_inAct_2,
  input  [15:0] io_inAct_3,
  input  [15:0] io_inAct_4,
  input  [15:0] io_inAct_5,
  input  [15:0] io_inAct_6,
  input  [15:0] io_inAct_7,
  input  [15:0] io_inAct_8,
  input  [15:0] io_inAct_9,
  input  [15:0] io_inAct_10,
  input  [15:0] io_inAct_11,
  input  [15:0] io_inAct_12,
  input  [15:0] io_inAct_13,
  input  [15:0] io_inAct_14,
  input  [15:0] io_inAct_15,
  input  [15:0] io_inAct_16,
  input  [15:0] io_inAct_17,
  input  [15:0] io_inAct_18,
  input  [15:0] io_inAct_19,
  input  [15:0] io_inWeight_0,
  input  [15:0] io_inWeight_1,
  input  [15:0] io_inWeight_2,
  input  [15:0] io_inWeight_3,
  input  [15:0] io_inWeight_4,
  input  [15:0] io_inWeight_5,
  input  [15:0] io_inWeight_6,
  input  [15:0] io_inWeight_7,
  input  [15:0] io_inWeight_8,
  input  [15:0] io_inWeight_9,
  output [39:0] io_outSum_0,
  output [39:0] io_outSum_1,
  output [39:0] io_outSum_2,
  output [39:0] io_outSum_3,
  output [39:0] io_outSum_4,
  output [39:0] io_outSum_5,
  output [39:0] io_outSum_6,
  output [39:0] io_outSum_7,
  output [39:0] io_outSum_8,
  output [39:0] io_outSum_9,
  input         io_inwtValid
);
  wire  PEs_0_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_10_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_10_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_10_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_10_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_11_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_11_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_11_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_11_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_12_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_12_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_12_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_12_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_13_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_13_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_13_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_13_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_14_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_14_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_14_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_14_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_15_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_15_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_15_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_15_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_16_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_16_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_16_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_16_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_17_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_17_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_17_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_17_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_18_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_18_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_18_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_18_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_19_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_19_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_19_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_19_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  reg  validReg; // @[SystolicArray.scala 22:25]
  PE PEs_0_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_0_clock),
    .io_inAct(PEs_0_0_io_inAct),
    .io_inWtPS(PEs_0_0_io_inWtPS),
    .io_outWtPS(PEs_0_0_io_outWtPS),
    .io_outAct(PEs_0_0_io_outAct),
    .io_inwtValid(PEs_0_0_io_inwtValid)
  );
  PE PEs_0_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_1_clock),
    .io_inAct(PEs_0_1_io_inAct),
    .io_inWtPS(PEs_0_1_io_inWtPS),
    .io_outWtPS(PEs_0_1_io_outWtPS),
    .io_outAct(PEs_0_1_io_outAct),
    .io_inwtValid(PEs_0_1_io_inwtValid)
  );
  PE PEs_0_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_2_clock),
    .io_inAct(PEs_0_2_io_inAct),
    .io_inWtPS(PEs_0_2_io_inWtPS),
    .io_outWtPS(PEs_0_2_io_outWtPS),
    .io_outAct(PEs_0_2_io_outAct),
    .io_inwtValid(PEs_0_2_io_inwtValid)
  );
  PE PEs_0_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_3_clock),
    .io_inAct(PEs_0_3_io_inAct),
    .io_inWtPS(PEs_0_3_io_inWtPS),
    .io_outWtPS(PEs_0_3_io_outWtPS),
    .io_outAct(PEs_0_3_io_outAct),
    .io_inwtValid(PEs_0_3_io_inwtValid)
  );
  PE PEs_0_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_4_clock),
    .io_inAct(PEs_0_4_io_inAct),
    .io_inWtPS(PEs_0_4_io_inWtPS),
    .io_outWtPS(PEs_0_4_io_outWtPS),
    .io_outAct(PEs_0_4_io_outAct),
    .io_inwtValid(PEs_0_4_io_inwtValid)
  );
  PE PEs_0_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_5_clock),
    .io_inAct(PEs_0_5_io_inAct),
    .io_inWtPS(PEs_0_5_io_inWtPS),
    .io_outWtPS(PEs_0_5_io_outWtPS),
    .io_outAct(PEs_0_5_io_outAct),
    .io_inwtValid(PEs_0_5_io_inwtValid)
  );
  PE PEs_0_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_6_clock),
    .io_inAct(PEs_0_6_io_inAct),
    .io_inWtPS(PEs_0_6_io_inWtPS),
    .io_outWtPS(PEs_0_6_io_outWtPS),
    .io_outAct(PEs_0_6_io_outAct),
    .io_inwtValid(PEs_0_6_io_inwtValid)
  );
  PE PEs_0_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_7_clock),
    .io_inAct(PEs_0_7_io_inAct),
    .io_inWtPS(PEs_0_7_io_inWtPS),
    .io_outWtPS(PEs_0_7_io_outWtPS),
    .io_outAct(PEs_0_7_io_outAct),
    .io_inwtValid(PEs_0_7_io_inwtValid)
  );
  PE PEs_0_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_8_clock),
    .io_inAct(PEs_0_8_io_inAct),
    .io_inWtPS(PEs_0_8_io_inWtPS),
    .io_outWtPS(PEs_0_8_io_outWtPS),
    .io_outAct(PEs_0_8_io_outAct),
    .io_inwtValid(PEs_0_8_io_inwtValid)
  );
  PE PEs_0_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_9_clock),
    .io_inAct(PEs_0_9_io_inAct),
    .io_inWtPS(PEs_0_9_io_inWtPS),
    .io_outWtPS(PEs_0_9_io_outWtPS),
    .io_outAct(PEs_0_9_io_outAct),
    .io_inwtValid(PEs_0_9_io_inwtValid)
  );
  PE PEs_1_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_0_clock),
    .io_inAct(PEs_1_0_io_inAct),
    .io_inWtPS(PEs_1_0_io_inWtPS),
    .io_outWtPS(PEs_1_0_io_outWtPS),
    .io_outAct(PEs_1_0_io_outAct),
    .io_inwtValid(PEs_1_0_io_inwtValid)
  );
  PE PEs_1_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_1_clock),
    .io_inAct(PEs_1_1_io_inAct),
    .io_inWtPS(PEs_1_1_io_inWtPS),
    .io_outWtPS(PEs_1_1_io_outWtPS),
    .io_outAct(PEs_1_1_io_outAct),
    .io_inwtValid(PEs_1_1_io_inwtValid)
  );
  PE PEs_1_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_2_clock),
    .io_inAct(PEs_1_2_io_inAct),
    .io_inWtPS(PEs_1_2_io_inWtPS),
    .io_outWtPS(PEs_1_2_io_outWtPS),
    .io_outAct(PEs_1_2_io_outAct),
    .io_inwtValid(PEs_1_2_io_inwtValid)
  );
  PE PEs_1_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_3_clock),
    .io_inAct(PEs_1_3_io_inAct),
    .io_inWtPS(PEs_1_3_io_inWtPS),
    .io_outWtPS(PEs_1_3_io_outWtPS),
    .io_outAct(PEs_1_3_io_outAct),
    .io_inwtValid(PEs_1_3_io_inwtValid)
  );
  PE PEs_1_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_4_clock),
    .io_inAct(PEs_1_4_io_inAct),
    .io_inWtPS(PEs_1_4_io_inWtPS),
    .io_outWtPS(PEs_1_4_io_outWtPS),
    .io_outAct(PEs_1_4_io_outAct),
    .io_inwtValid(PEs_1_4_io_inwtValid)
  );
  PE PEs_1_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_5_clock),
    .io_inAct(PEs_1_5_io_inAct),
    .io_inWtPS(PEs_1_5_io_inWtPS),
    .io_outWtPS(PEs_1_5_io_outWtPS),
    .io_outAct(PEs_1_5_io_outAct),
    .io_inwtValid(PEs_1_5_io_inwtValid)
  );
  PE PEs_1_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_6_clock),
    .io_inAct(PEs_1_6_io_inAct),
    .io_inWtPS(PEs_1_6_io_inWtPS),
    .io_outWtPS(PEs_1_6_io_outWtPS),
    .io_outAct(PEs_1_6_io_outAct),
    .io_inwtValid(PEs_1_6_io_inwtValid)
  );
  PE PEs_1_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_7_clock),
    .io_inAct(PEs_1_7_io_inAct),
    .io_inWtPS(PEs_1_7_io_inWtPS),
    .io_outWtPS(PEs_1_7_io_outWtPS),
    .io_outAct(PEs_1_7_io_outAct),
    .io_inwtValid(PEs_1_7_io_inwtValid)
  );
  PE PEs_1_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_8_clock),
    .io_inAct(PEs_1_8_io_inAct),
    .io_inWtPS(PEs_1_8_io_inWtPS),
    .io_outWtPS(PEs_1_8_io_outWtPS),
    .io_outAct(PEs_1_8_io_outAct),
    .io_inwtValid(PEs_1_8_io_inwtValid)
  );
  PE PEs_1_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_9_clock),
    .io_inAct(PEs_1_9_io_inAct),
    .io_inWtPS(PEs_1_9_io_inWtPS),
    .io_outWtPS(PEs_1_9_io_outWtPS),
    .io_outAct(PEs_1_9_io_outAct),
    .io_inwtValid(PEs_1_9_io_inwtValid)
  );
  PE PEs_2_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_0_clock),
    .io_inAct(PEs_2_0_io_inAct),
    .io_inWtPS(PEs_2_0_io_inWtPS),
    .io_outWtPS(PEs_2_0_io_outWtPS),
    .io_outAct(PEs_2_0_io_outAct),
    .io_inwtValid(PEs_2_0_io_inwtValid)
  );
  PE PEs_2_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_1_clock),
    .io_inAct(PEs_2_1_io_inAct),
    .io_inWtPS(PEs_2_1_io_inWtPS),
    .io_outWtPS(PEs_2_1_io_outWtPS),
    .io_outAct(PEs_2_1_io_outAct),
    .io_inwtValid(PEs_2_1_io_inwtValid)
  );
  PE PEs_2_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_2_clock),
    .io_inAct(PEs_2_2_io_inAct),
    .io_inWtPS(PEs_2_2_io_inWtPS),
    .io_outWtPS(PEs_2_2_io_outWtPS),
    .io_outAct(PEs_2_2_io_outAct),
    .io_inwtValid(PEs_2_2_io_inwtValid)
  );
  PE PEs_2_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_3_clock),
    .io_inAct(PEs_2_3_io_inAct),
    .io_inWtPS(PEs_2_3_io_inWtPS),
    .io_outWtPS(PEs_2_3_io_outWtPS),
    .io_outAct(PEs_2_3_io_outAct),
    .io_inwtValid(PEs_2_3_io_inwtValid)
  );
  PE PEs_2_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_4_clock),
    .io_inAct(PEs_2_4_io_inAct),
    .io_inWtPS(PEs_2_4_io_inWtPS),
    .io_outWtPS(PEs_2_4_io_outWtPS),
    .io_outAct(PEs_2_4_io_outAct),
    .io_inwtValid(PEs_2_4_io_inwtValid)
  );
  PE PEs_2_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_5_clock),
    .io_inAct(PEs_2_5_io_inAct),
    .io_inWtPS(PEs_2_5_io_inWtPS),
    .io_outWtPS(PEs_2_5_io_outWtPS),
    .io_outAct(PEs_2_5_io_outAct),
    .io_inwtValid(PEs_2_5_io_inwtValid)
  );
  PE PEs_2_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_6_clock),
    .io_inAct(PEs_2_6_io_inAct),
    .io_inWtPS(PEs_2_6_io_inWtPS),
    .io_outWtPS(PEs_2_6_io_outWtPS),
    .io_outAct(PEs_2_6_io_outAct),
    .io_inwtValid(PEs_2_6_io_inwtValid)
  );
  PE PEs_2_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_7_clock),
    .io_inAct(PEs_2_7_io_inAct),
    .io_inWtPS(PEs_2_7_io_inWtPS),
    .io_outWtPS(PEs_2_7_io_outWtPS),
    .io_outAct(PEs_2_7_io_outAct),
    .io_inwtValid(PEs_2_7_io_inwtValid)
  );
  PE PEs_2_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_8_clock),
    .io_inAct(PEs_2_8_io_inAct),
    .io_inWtPS(PEs_2_8_io_inWtPS),
    .io_outWtPS(PEs_2_8_io_outWtPS),
    .io_outAct(PEs_2_8_io_outAct),
    .io_inwtValid(PEs_2_8_io_inwtValid)
  );
  PE PEs_2_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_9_clock),
    .io_inAct(PEs_2_9_io_inAct),
    .io_inWtPS(PEs_2_9_io_inWtPS),
    .io_outWtPS(PEs_2_9_io_outWtPS),
    .io_outAct(PEs_2_9_io_outAct),
    .io_inwtValid(PEs_2_9_io_inwtValid)
  );
  PE PEs_3_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_0_clock),
    .io_inAct(PEs_3_0_io_inAct),
    .io_inWtPS(PEs_3_0_io_inWtPS),
    .io_outWtPS(PEs_3_0_io_outWtPS),
    .io_outAct(PEs_3_0_io_outAct),
    .io_inwtValid(PEs_3_0_io_inwtValid)
  );
  PE PEs_3_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_1_clock),
    .io_inAct(PEs_3_1_io_inAct),
    .io_inWtPS(PEs_3_1_io_inWtPS),
    .io_outWtPS(PEs_3_1_io_outWtPS),
    .io_outAct(PEs_3_1_io_outAct),
    .io_inwtValid(PEs_3_1_io_inwtValid)
  );
  PE PEs_3_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_2_clock),
    .io_inAct(PEs_3_2_io_inAct),
    .io_inWtPS(PEs_3_2_io_inWtPS),
    .io_outWtPS(PEs_3_2_io_outWtPS),
    .io_outAct(PEs_3_2_io_outAct),
    .io_inwtValid(PEs_3_2_io_inwtValid)
  );
  PE PEs_3_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_3_clock),
    .io_inAct(PEs_3_3_io_inAct),
    .io_inWtPS(PEs_3_3_io_inWtPS),
    .io_outWtPS(PEs_3_3_io_outWtPS),
    .io_outAct(PEs_3_3_io_outAct),
    .io_inwtValid(PEs_3_3_io_inwtValid)
  );
  PE PEs_3_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_4_clock),
    .io_inAct(PEs_3_4_io_inAct),
    .io_inWtPS(PEs_3_4_io_inWtPS),
    .io_outWtPS(PEs_3_4_io_outWtPS),
    .io_outAct(PEs_3_4_io_outAct),
    .io_inwtValid(PEs_3_4_io_inwtValid)
  );
  PE PEs_3_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_5_clock),
    .io_inAct(PEs_3_5_io_inAct),
    .io_inWtPS(PEs_3_5_io_inWtPS),
    .io_outWtPS(PEs_3_5_io_outWtPS),
    .io_outAct(PEs_3_5_io_outAct),
    .io_inwtValid(PEs_3_5_io_inwtValid)
  );
  PE PEs_3_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_6_clock),
    .io_inAct(PEs_3_6_io_inAct),
    .io_inWtPS(PEs_3_6_io_inWtPS),
    .io_outWtPS(PEs_3_6_io_outWtPS),
    .io_outAct(PEs_3_6_io_outAct),
    .io_inwtValid(PEs_3_6_io_inwtValid)
  );
  PE PEs_3_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_7_clock),
    .io_inAct(PEs_3_7_io_inAct),
    .io_inWtPS(PEs_3_7_io_inWtPS),
    .io_outWtPS(PEs_3_7_io_outWtPS),
    .io_outAct(PEs_3_7_io_outAct),
    .io_inwtValid(PEs_3_7_io_inwtValid)
  );
  PE PEs_3_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_8_clock),
    .io_inAct(PEs_3_8_io_inAct),
    .io_inWtPS(PEs_3_8_io_inWtPS),
    .io_outWtPS(PEs_3_8_io_outWtPS),
    .io_outAct(PEs_3_8_io_outAct),
    .io_inwtValid(PEs_3_8_io_inwtValid)
  );
  PE PEs_3_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_9_clock),
    .io_inAct(PEs_3_9_io_inAct),
    .io_inWtPS(PEs_3_9_io_inWtPS),
    .io_outWtPS(PEs_3_9_io_outWtPS),
    .io_outAct(PEs_3_9_io_outAct),
    .io_inwtValid(PEs_3_9_io_inwtValid)
  );
  PE PEs_4_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_0_clock),
    .io_inAct(PEs_4_0_io_inAct),
    .io_inWtPS(PEs_4_0_io_inWtPS),
    .io_outWtPS(PEs_4_0_io_outWtPS),
    .io_outAct(PEs_4_0_io_outAct),
    .io_inwtValid(PEs_4_0_io_inwtValid)
  );
  PE PEs_4_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_1_clock),
    .io_inAct(PEs_4_1_io_inAct),
    .io_inWtPS(PEs_4_1_io_inWtPS),
    .io_outWtPS(PEs_4_1_io_outWtPS),
    .io_outAct(PEs_4_1_io_outAct),
    .io_inwtValid(PEs_4_1_io_inwtValid)
  );
  PE PEs_4_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_2_clock),
    .io_inAct(PEs_4_2_io_inAct),
    .io_inWtPS(PEs_4_2_io_inWtPS),
    .io_outWtPS(PEs_4_2_io_outWtPS),
    .io_outAct(PEs_4_2_io_outAct),
    .io_inwtValid(PEs_4_2_io_inwtValid)
  );
  PE PEs_4_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_3_clock),
    .io_inAct(PEs_4_3_io_inAct),
    .io_inWtPS(PEs_4_3_io_inWtPS),
    .io_outWtPS(PEs_4_3_io_outWtPS),
    .io_outAct(PEs_4_3_io_outAct),
    .io_inwtValid(PEs_4_3_io_inwtValid)
  );
  PE PEs_4_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_4_clock),
    .io_inAct(PEs_4_4_io_inAct),
    .io_inWtPS(PEs_4_4_io_inWtPS),
    .io_outWtPS(PEs_4_4_io_outWtPS),
    .io_outAct(PEs_4_4_io_outAct),
    .io_inwtValid(PEs_4_4_io_inwtValid)
  );
  PE PEs_4_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_5_clock),
    .io_inAct(PEs_4_5_io_inAct),
    .io_inWtPS(PEs_4_5_io_inWtPS),
    .io_outWtPS(PEs_4_5_io_outWtPS),
    .io_outAct(PEs_4_5_io_outAct),
    .io_inwtValid(PEs_4_5_io_inwtValid)
  );
  PE PEs_4_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_6_clock),
    .io_inAct(PEs_4_6_io_inAct),
    .io_inWtPS(PEs_4_6_io_inWtPS),
    .io_outWtPS(PEs_4_6_io_outWtPS),
    .io_outAct(PEs_4_6_io_outAct),
    .io_inwtValid(PEs_4_6_io_inwtValid)
  );
  PE PEs_4_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_7_clock),
    .io_inAct(PEs_4_7_io_inAct),
    .io_inWtPS(PEs_4_7_io_inWtPS),
    .io_outWtPS(PEs_4_7_io_outWtPS),
    .io_outAct(PEs_4_7_io_outAct),
    .io_inwtValid(PEs_4_7_io_inwtValid)
  );
  PE PEs_4_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_8_clock),
    .io_inAct(PEs_4_8_io_inAct),
    .io_inWtPS(PEs_4_8_io_inWtPS),
    .io_outWtPS(PEs_4_8_io_outWtPS),
    .io_outAct(PEs_4_8_io_outAct),
    .io_inwtValid(PEs_4_8_io_inwtValid)
  );
  PE PEs_4_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_9_clock),
    .io_inAct(PEs_4_9_io_inAct),
    .io_inWtPS(PEs_4_9_io_inWtPS),
    .io_outWtPS(PEs_4_9_io_outWtPS),
    .io_outAct(PEs_4_9_io_outAct),
    .io_inwtValid(PEs_4_9_io_inwtValid)
  );
  PE PEs_5_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_0_clock),
    .io_inAct(PEs_5_0_io_inAct),
    .io_inWtPS(PEs_5_0_io_inWtPS),
    .io_outWtPS(PEs_5_0_io_outWtPS),
    .io_outAct(PEs_5_0_io_outAct),
    .io_inwtValid(PEs_5_0_io_inwtValid)
  );
  PE PEs_5_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_1_clock),
    .io_inAct(PEs_5_1_io_inAct),
    .io_inWtPS(PEs_5_1_io_inWtPS),
    .io_outWtPS(PEs_5_1_io_outWtPS),
    .io_outAct(PEs_5_1_io_outAct),
    .io_inwtValid(PEs_5_1_io_inwtValid)
  );
  PE PEs_5_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_2_clock),
    .io_inAct(PEs_5_2_io_inAct),
    .io_inWtPS(PEs_5_2_io_inWtPS),
    .io_outWtPS(PEs_5_2_io_outWtPS),
    .io_outAct(PEs_5_2_io_outAct),
    .io_inwtValid(PEs_5_2_io_inwtValid)
  );
  PE PEs_5_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_3_clock),
    .io_inAct(PEs_5_3_io_inAct),
    .io_inWtPS(PEs_5_3_io_inWtPS),
    .io_outWtPS(PEs_5_3_io_outWtPS),
    .io_outAct(PEs_5_3_io_outAct),
    .io_inwtValid(PEs_5_3_io_inwtValid)
  );
  PE PEs_5_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_4_clock),
    .io_inAct(PEs_5_4_io_inAct),
    .io_inWtPS(PEs_5_4_io_inWtPS),
    .io_outWtPS(PEs_5_4_io_outWtPS),
    .io_outAct(PEs_5_4_io_outAct),
    .io_inwtValid(PEs_5_4_io_inwtValid)
  );
  PE PEs_5_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_5_clock),
    .io_inAct(PEs_5_5_io_inAct),
    .io_inWtPS(PEs_5_5_io_inWtPS),
    .io_outWtPS(PEs_5_5_io_outWtPS),
    .io_outAct(PEs_5_5_io_outAct),
    .io_inwtValid(PEs_5_5_io_inwtValid)
  );
  PE PEs_5_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_6_clock),
    .io_inAct(PEs_5_6_io_inAct),
    .io_inWtPS(PEs_5_6_io_inWtPS),
    .io_outWtPS(PEs_5_6_io_outWtPS),
    .io_outAct(PEs_5_6_io_outAct),
    .io_inwtValid(PEs_5_6_io_inwtValid)
  );
  PE PEs_5_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_7_clock),
    .io_inAct(PEs_5_7_io_inAct),
    .io_inWtPS(PEs_5_7_io_inWtPS),
    .io_outWtPS(PEs_5_7_io_outWtPS),
    .io_outAct(PEs_5_7_io_outAct),
    .io_inwtValid(PEs_5_7_io_inwtValid)
  );
  PE PEs_5_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_8_clock),
    .io_inAct(PEs_5_8_io_inAct),
    .io_inWtPS(PEs_5_8_io_inWtPS),
    .io_outWtPS(PEs_5_8_io_outWtPS),
    .io_outAct(PEs_5_8_io_outAct),
    .io_inwtValid(PEs_5_8_io_inwtValid)
  );
  PE PEs_5_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_9_clock),
    .io_inAct(PEs_5_9_io_inAct),
    .io_inWtPS(PEs_5_9_io_inWtPS),
    .io_outWtPS(PEs_5_9_io_outWtPS),
    .io_outAct(PEs_5_9_io_outAct),
    .io_inwtValid(PEs_5_9_io_inwtValid)
  );
  PE PEs_6_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_0_clock),
    .io_inAct(PEs_6_0_io_inAct),
    .io_inWtPS(PEs_6_0_io_inWtPS),
    .io_outWtPS(PEs_6_0_io_outWtPS),
    .io_outAct(PEs_6_0_io_outAct),
    .io_inwtValid(PEs_6_0_io_inwtValid)
  );
  PE PEs_6_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_1_clock),
    .io_inAct(PEs_6_1_io_inAct),
    .io_inWtPS(PEs_6_1_io_inWtPS),
    .io_outWtPS(PEs_6_1_io_outWtPS),
    .io_outAct(PEs_6_1_io_outAct),
    .io_inwtValid(PEs_6_1_io_inwtValid)
  );
  PE PEs_6_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_2_clock),
    .io_inAct(PEs_6_2_io_inAct),
    .io_inWtPS(PEs_6_2_io_inWtPS),
    .io_outWtPS(PEs_6_2_io_outWtPS),
    .io_outAct(PEs_6_2_io_outAct),
    .io_inwtValid(PEs_6_2_io_inwtValid)
  );
  PE PEs_6_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_3_clock),
    .io_inAct(PEs_6_3_io_inAct),
    .io_inWtPS(PEs_6_3_io_inWtPS),
    .io_outWtPS(PEs_6_3_io_outWtPS),
    .io_outAct(PEs_6_3_io_outAct),
    .io_inwtValid(PEs_6_3_io_inwtValid)
  );
  PE PEs_6_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_4_clock),
    .io_inAct(PEs_6_4_io_inAct),
    .io_inWtPS(PEs_6_4_io_inWtPS),
    .io_outWtPS(PEs_6_4_io_outWtPS),
    .io_outAct(PEs_6_4_io_outAct),
    .io_inwtValid(PEs_6_4_io_inwtValid)
  );
  PE PEs_6_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_5_clock),
    .io_inAct(PEs_6_5_io_inAct),
    .io_inWtPS(PEs_6_5_io_inWtPS),
    .io_outWtPS(PEs_6_5_io_outWtPS),
    .io_outAct(PEs_6_5_io_outAct),
    .io_inwtValid(PEs_6_5_io_inwtValid)
  );
  PE PEs_6_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_6_clock),
    .io_inAct(PEs_6_6_io_inAct),
    .io_inWtPS(PEs_6_6_io_inWtPS),
    .io_outWtPS(PEs_6_6_io_outWtPS),
    .io_outAct(PEs_6_6_io_outAct),
    .io_inwtValid(PEs_6_6_io_inwtValid)
  );
  PE PEs_6_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_7_clock),
    .io_inAct(PEs_6_7_io_inAct),
    .io_inWtPS(PEs_6_7_io_inWtPS),
    .io_outWtPS(PEs_6_7_io_outWtPS),
    .io_outAct(PEs_6_7_io_outAct),
    .io_inwtValid(PEs_6_7_io_inwtValid)
  );
  PE PEs_6_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_8_clock),
    .io_inAct(PEs_6_8_io_inAct),
    .io_inWtPS(PEs_6_8_io_inWtPS),
    .io_outWtPS(PEs_6_8_io_outWtPS),
    .io_outAct(PEs_6_8_io_outAct),
    .io_inwtValid(PEs_6_8_io_inwtValid)
  );
  PE PEs_6_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_9_clock),
    .io_inAct(PEs_6_9_io_inAct),
    .io_inWtPS(PEs_6_9_io_inWtPS),
    .io_outWtPS(PEs_6_9_io_outWtPS),
    .io_outAct(PEs_6_9_io_outAct),
    .io_inwtValid(PEs_6_9_io_inwtValid)
  );
  PE PEs_7_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_0_clock),
    .io_inAct(PEs_7_0_io_inAct),
    .io_inWtPS(PEs_7_0_io_inWtPS),
    .io_outWtPS(PEs_7_0_io_outWtPS),
    .io_outAct(PEs_7_0_io_outAct),
    .io_inwtValid(PEs_7_0_io_inwtValid)
  );
  PE PEs_7_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_1_clock),
    .io_inAct(PEs_7_1_io_inAct),
    .io_inWtPS(PEs_7_1_io_inWtPS),
    .io_outWtPS(PEs_7_1_io_outWtPS),
    .io_outAct(PEs_7_1_io_outAct),
    .io_inwtValid(PEs_7_1_io_inwtValid)
  );
  PE PEs_7_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_2_clock),
    .io_inAct(PEs_7_2_io_inAct),
    .io_inWtPS(PEs_7_2_io_inWtPS),
    .io_outWtPS(PEs_7_2_io_outWtPS),
    .io_outAct(PEs_7_2_io_outAct),
    .io_inwtValid(PEs_7_2_io_inwtValid)
  );
  PE PEs_7_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_3_clock),
    .io_inAct(PEs_7_3_io_inAct),
    .io_inWtPS(PEs_7_3_io_inWtPS),
    .io_outWtPS(PEs_7_3_io_outWtPS),
    .io_outAct(PEs_7_3_io_outAct),
    .io_inwtValid(PEs_7_3_io_inwtValid)
  );
  PE PEs_7_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_4_clock),
    .io_inAct(PEs_7_4_io_inAct),
    .io_inWtPS(PEs_7_4_io_inWtPS),
    .io_outWtPS(PEs_7_4_io_outWtPS),
    .io_outAct(PEs_7_4_io_outAct),
    .io_inwtValid(PEs_7_4_io_inwtValid)
  );
  PE PEs_7_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_5_clock),
    .io_inAct(PEs_7_5_io_inAct),
    .io_inWtPS(PEs_7_5_io_inWtPS),
    .io_outWtPS(PEs_7_5_io_outWtPS),
    .io_outAct(PEs_7_5_io_outAct),
    .io_inwtValid(PEs_7_5_io_inwtValid)
  );
  PE PEs_7_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_6_clock),
    .io_inAct(PEs_7_6_io_inAct),
    .io_inWtPS(PEs_7_6_io_inWtPS),
    .io_outWtPS(PEs_7_6_io_outWtPS),
    .io_outAct(PEs_7_6_io_outAct),
    .io_inwtValid(PEs_7_6_io_inwtValid)
  );
  PE PEs_7_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_7_clock),
    .io_inAct(PEs_7_7_io_inAct),
    .io_inWtPS(PEs_7_7_io_inWtPS),
    .io_outWtPS(PEs_7_7_io_outWtPS),
    .io_outAct(PEs_7_7_io_outAct),
    .io_inwtValid(PEs_7_7_io_inwtValid)
  );
  PE PEs_7_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_8_clock),
    .io_inAct(PEs_7_8_io_inAct),
    .io_inWtPS(PEs_7_8_io_inWtPS),
    .io_outWtPS(PEs_7_8_io_outWtPS),
    .io_outAct(PEs_7_8_io_outAct),
    .io_inwtValid(PEs_7_8_io_inwtValid)
  );
  PE PEs_7_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_9_clock),
    .io_inAct(PEs_7_9_io_inAct),
    .io_inWtPS(PEs_7_9_io_inWtPS),
    .io_outWtPS(PEs_7_9_io_outWtPS),
    .io_outAct(PEs_7_9_io_outAct),
    .io_inwtValid(PEs_7_9_io_inwtValid)
  );
  PE PEs_8_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_0_clock),
    .io_inAct(PEs_8_0_io_inAct),
    .io_inWtPS(PEs_8_0_io_inWtPS),
    .io_outWtPS(PEs_8_0_io_outWtPS),
    .io_outAct(PEs_8_0_io_outAct),
    .io_inwtValid(PEs_8_0_io_inwtValid)
  );
  PE PEs_8_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_1_clock),
    .io_inAct(PEs_8_1_io_inAct),
    .io_inWtPS(PEs_8_1_io_inWtPS),
    .io_outWtPS(PEs_8_1_io_outWtPS),
    .io_outAct(PEs_8_1_io_outAct),
    .io_inwtValid(PEs_8_1_io_inwtValid)
  );
  PE PEs_8_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_2_clock),
    .io_inAct(PEs_8_2_io_inAct),
    .io_inWtPS(PEs_8_2_io_inWtPS),
    .io_outWtPS(PEs_8_2_io_outWtPS),
    .io_outAct(PEs_8_2_io_outAct),
    .io_inwtValid(PEs_8_2_io_inwtValid)
  );
  PE PEs_8_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_3_clock),
    .io_inAct(PEs_8_3_io_inAct),
    .io_inWtPS(PEs_8_3_io_inWtPS),
    .io_outWtPS(PEs_8_3_io_outWtPS),
    .io_outAct(PEs_8_3_io_outAct),
    .io_inwtValid(PEs_8_3_io_inwtValid)
  );
  PE PEs_8_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_4_clock),
    .io_inAct(PEs_8_4_io_inAct),
    .io_inWtPS(PEs_8_4_io_inWtPS),
    .io_outWtPS(PEs_8_4_io_outWtPS),
    .io_outAct(PEs_8_4_io_outAct),
    .io_inwtValid(PEs_8_4_io_inwtValid)
  );
  PE PEs_8_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_5_clock),
    .io_inAct(PEs_8_5_io_inAct),
    .io_inWtPS(PEs_8_5_io_inWtPS),
    .io_outWtPS(PEs_8_5_io_outWtPS),
    .io_outAct(PEs_8_5_io_outAct),
    .io_inwtValid(PEs_8_5_io_inwtValid)
  );
  PE PEs_8_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_6_clock),
    .io_inAct(PEs_8_6_io_inAct),
    .io_inWtPS(PEs_8_6_io_inWtPS),
    .io_outWtPS(PEs_8_6_io_outWtPS),
    .io_outAct(PEs_8_6_io_outAct),
    .io_inwtValid(PEs_8_6_io_inwtValid)
  );
  PE PEs_8_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_7_clock),
    .io_inAct(PEs_8_7_io_inAct),
    .io_inWtPS(PEs_8_7_io_inWtPS),
    .io_outWtPS(PEs_8_7_io_outWtPS),
    .io_outAct(PEs_8_7_io_outAct),
    .io_inwtValid(PEs_8_7_io_inwtValid)
  );
  PE PEs_8_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_8_clock),
    .io_inAct(PEs_8_8_io_inAct),
    .io_inWtPS(PEs_8_8_io_inWtPS),
    .io_outWtPS(PEs_8_8_io_outWtPS),
    .io_outAct(PEs_8_8_io_outAct),
    .io_inwtValid(PEs_8_8_io_inwtValid)
  );
  PE PEs_8_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_9_clock),
    .io_inAct(PEs_8_9_io_inAct),
    .io_inWtPS(PEs_8_9_io_inWtPS),
    .io_outWtPS(PEs_8_9_io_outWtPS),
    .io_outAct(PEs_8_9_io_outAct),
    .io_inwtValid(PEs_8_9_io_inwtValid)
  );
  PE PEs_9_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_0_clock),
    .io_inAct(PEs_9_0_io_inAct),
    .io_inWtPS(PEs_9_0_io_inWtPS),
    .io_outWtPS(PEs_9_0_io_outWtPS),
    .io_outAct(PEs_9_0_io_outAct),
    .io_inwtValid(PEs_9_0_io_inwtValid)
  );
  PE PEs_9_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_1_clock),
    .io_inAct(PEs_9_1_io_inAct),
    .io_inWtPS(PEs_9_1_io_inWtPS),
    .io_outWtPS(PEs_9_1_io_outWtPS),
    .io_outAct(PEs_9_1_io_outAct),
    .io_inwtValid(PEs_9_1_io_inwtValid)
  );
  PE PEs_9_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_2_clock),
    .io_inAct(PEs_9_2_io_inAct),
    .io_inWtPS(PEs_9_2_io_inWtPS),
    .io_outWtPS(PEs_9_2_io_outWtPS),
    .io_outAct(PEs_9_2_io_outAct),
    .io_inwtValid(PEs_9_2_io_inwtValid)
  );
  PE PEs_9_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_3_clock),
    .io_inAct(PEs_9_3_io_inAct),
    .io_inWtPS(PEs_9_3_io_inWtPS),
    .io_outWtPS(PEs_9_3_io_outWtPS),
    .io_outAct(PEs_9_3_io_outAct),
    .io_inwtValid(PEs_9_3_io_inwtValid)
  );
  PE PEs_9_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_4_clock),
    .io_inAct(PEs_9_4_io_inAct),
    .io_inWtPS(PEs_9_4_io_inWtPS),
    .io_outWtPS(PEs_9_4_io_outWtPS),
    .io_outAct(PEs_9_4_io_outAct),
    .io_inwtValid(PEs_9_4_io_inwtValid)
  );
  PE PEs_9_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_5_clock),
    .io_inAct(PEs_9_5_io_inAct),
    .io_inWtPS(PEs_9_5_io_inWtPS),
    .io_outWtPS(PEs_9_5_io_outWtPS),
    .io_outAct(PEs_9_5_io_outAct),
    .io_inwtValid(PEs_9_5_io_inwtValid)
  );
  PE PEs_9_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_6_clock),
    .io_inAct(PEs_9_6_io_inAct),
    .io_inWtPS(PEs_9_6_io_inWtPS),
    .io_outWtPS(PEs_9_6_io_outWtPS),
    .io_outAct(PEs_9_6_io_outAct),
    .io_inwtValid(PEs_9_6_io_inwtValid)
  );
  PE PEs_9_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_7_clock),
    .io_inAct(PEs_9_7_io_inAct),
    .io_inWtPS(PEs_9_7_io_inWtPS),
    .io_outWtPS(PEs_9_7_io_outWtPS),
    .io_outAct(PEs_9_7_io_outAct),
    .io_inwtValid(PEs_9_7_io_inwtValid)
  );
  PE PEs_9_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_8_clock),
    .io_inAct(PEs_9_8_io_inAct),
    .io_inWtPS(PEs_9_8_io_inWtPS),
    .io_outWtPS(PEs_9_8_io_outWtPS),
    .io_outAct(PEs_9_8_io_outAct),
    .io_inwtValid(PEs_9_8_io_inwtValid)
  );
  PE PEs_9_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_9_clock),
    .io_inAct(PEs_9_9_io_inAct),
    .io_inWtPS(PEs_9_9_io_inWtPS),
    .io_outWtPS(PEs_9_9_io_outWtPS),
    .io_outAct(PEs_9_9_io_outAct),
    .io_inwtValid(PEs_9_9_io_inwtValid)
  );
  PE PEs_10_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_0_clock),
    .io_inAct(PEs_10_0_io_inAct),
    .io_inWtPS(PEs_10_0_io_inWtPS),
    .io_outWtPS(PEs_10_0_io_outWtPS),
    .io_outAct(PEs_10_0_io_outAct),
    .io_inwtValid(PEs_10_0_io_inwtValid)
  );
  PE PEs_10_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_1_clock),
    .io_inAct(PEs_10_1_io_inAct),
    .io_inWtPS(PEs_10_1_io_inWtPS),
    .io_outWtPS(PEs_10_1_io_outWtPS),
    .io_outAct(PEs_10_1_io_outAct),
    .io_inwtValid(PEs_10_1_io_inwtValid)
  );
  PE PEs_10_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_2_clock),
    .io_inAct(PEs_10_2_io_inAct),
    .io_inWtPS(PEs_10_2_io_inWtPS),
    .io_outWtPS(PEs_10_2_io_outWtPS),
    .io_outAct(PEs_10_2_io_outAct),
    .io_inwtValid(PEs_10_2_io_inwtValid)
  );
  PE PEs_10_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_3_clock),
    .io_inAct(PEs_10_3_io_inAct),
    .io_inWtPS(PEs_10_3_io_inWtPS),
    .io_outWtPS(PEs_10_3_io_outWtPS),
    .io_outAct(PEs_10_3_io_outAct),
    .io_inwtValid(PEs_10_3_io_inwtValid)
  );
  PE PEs_10_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_4_clock),
    .io_inAct(PEs_10_4_io_inAct),
    .io_inWtPS(PEs_10_4_io_inWtPS),
    .io_outWtPS(PEs_10_4_io_outWtPS),
    .io_outAct(PEs_10_4_io_outAct),
    .io_inwtValid(PEs_10_4_io_inwtValid)
  );
  PE PEs_10_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_5_clock),
    .io_inAct(PEs_10_5_io_inAct),
    .io_inWtPS(PEs_10_5_io_inWtPS),
    .io_outWtPS(PEs_10_5_io_outWtPS),
    .io_outAct(PEs_10_5_io_outAct),
    .io_inwtValid(PEs_10_5_io_inwtValid)
  );
  PE PEs_10_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_6_clock),
    .io_inAct(PEs_10_6_io_inAct),
    .io_inWtPS(PEs_10_6_io_inWtPS),
    .io_outWtPS(PEs_10_6_io_outWtPS),
    .io_outAct(PEs_10_6_io_outAct),
    .io_inwtValid(PEs_10_6_io_inwtValid)
  );
  PE PEs_10_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_7_clock),
    .io_inAct(PEs_10_7_io_inAct),
    .io_inWtPS(PEs_10_7_io_inWtPS),
    .io_outWtPS(PEs_10_7_io_outWtPS),
    .io_outAct(PEs_10_7_io_outAct),
    .io_inwtValid(PEs_10_7_io_inwtValid)
  );
  PE PEs_10_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_8_clock),
    .io_inAct(PEs_10_8_io_inAct),
    .io_inWtPS(PEs_10_8_io_inWtPS),
    .io_outWtPS(PEs_10_8_io_outWtPS),
    .io_outAct(PEs_10_8_io_outAct),
    .io_inwtValid(PEs_10_8_io_inwtValid)
  );
  PE PEs_10_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_10_9_clock),
    .io_inAct(PEs_10_9_io_inAct),
    .io_inWtPS(PEs_10_9_io_inWtPS),
    .io_outWtPS(PEs_10_9_io_outWtPS),
    .io_outAct(PEs_10_9_io_outAct),
    .io_inwtValid(PEs_10_9_io_inwtValid)
  );
  PE PEs_11_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_0_clock),
    .io_inAct(PEs_11_0_io_inAct),
    .io_inWtPS(PEs_11_0_io_inWtPS),
    .io_outWtPS(PEs_11_0_io_outWtPS),
    .io_outAct(PEs_11_0_io_outAct),
    .io_inwtValid(PEs_11_0_io_inwtValid)
  );
  PE PEs_11_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_1_clock),
    .io_inAct(PEs_11_1_io_inAct),
    .io_inWtPS(PEs_11_1_io_inWtPS),
    .io_outWtPS(PEs_11_1_io_outWtPS),
    .io_outAct(PEs_11_1_io_outAct),
    .io_inwtValid(PEs_11_1_io_inwtValid)
  );
  PE PEs_11_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_2_clock),
    .io_inAct(PEs_11_2_io_inAct),
    .io_inWtPS(PEs_11_2_io_inWtPS),
    .io_outWtPS(PEs_11_2_io_outWtPS),
    .io_outAct(PEs_11_2_io_outAct),
    .io_inwtValid(PEs_11_2_io_inwtValid)
  );
  PE PEs_11_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_3_clock),
    .io_inAct(PEs_11_3_io_inAct),
    .io_inWtPS(PEs_11_3_io_inWtPS),
    .io_outWtPS(PEs_11_3_io_outWtPS),
    .io_outAct(PEs_11_3_io_outAct),
    .io_inwtValid(PEs_11_3_io_inwtValid)
  );
  PE PEs_11_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_4_clock),
    .io_inAct(PEs_11_4_io_inAct),
    .io_inWtPS(PEs_11_4_io_inWtPS),
    .io_outWtPS(PEs_11_4_io_outWtPS),
    .io_outAct(PEs_11_4_io_outAct),
    .io_inwtValid(PEs_11_4_io_inwtValid)
  );
  PE PEs_11_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_5_clock),
    .io_inAct(PEs_11_5_io_inAct),
    .io_inWtPS(PEs_11_5_io_inWtPS),
    .io_outWtPS(PEs_11_5_io_outWtPS),
    .io_outAct(PEs_11_5_io_outAct),
    .io_inwtValid(PEs_11_5_io_inwtValid)
  );
  PE PEs_11_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_6_clock),
    .io_inAct(PEs_11_6_io_inAct),
    .io_inWtPS(PEs_11_6_io_inWtPS),
    .io_outWtPS(PEs_11_6_io_outWtPS),
    .io_outAct(PEs_11_6_io_outAct),
    .io_inwtValid(PEs_11_6_io_inwtValid)
  );
  PE PEs_11_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_7_clock),
    .io_inAct(PEs_11_7_io_inAct),
    .io_inWtPS(PEs_11_7_io_inWtPS),
    .io_outWtPS(PEs_11_7_io_outWtPS),
    .io_outAct(PEs_11_7_io_outAct),
    .io_inwtValid(PEs_11_7_io_inwtValid)
  );
  PE PEs_11_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_8_clock),
    .io_inAct(PEs_11_8_io_inAct),
    .io_inWtPS(PEs_11_8_io_inWtPS),
    .io_outWtPS(PEs_11_8_io_outWtPS),
    .io_outAct(PEs_11_8_io_outAct),
    .io_inwtValid(PEs_11_8_io_inwtValid)
  );
  PE PEs_11_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_11_9_clock),
    .io_inAct(PEs_11_9_io_inAct),
    .io_inWtPS(PEs_11_9_io_inWtPS),
    .io_outWtPS(PEs_11_9_io_outWtPS),
    .io_outAct(PEs_11_9_io_outAct),
    .io_inwtValid(PEs_11_9_io_inwtValid)
  );
  PE PEs_12_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_0_clock),
    .io_inAct(PEs_12_0_io_inAct),
    .io_inWtPS(PEs_12_0_io_inWtPS),
    .io_outWtPS(PEs_12_0_io_outWtPS),
    .io_outAct(PEs_12_0_io_outAct),
    .io_inwtValid(PEs_12_0_io_inwtValid)
  );
  PE PEs_12_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_1_clock),
    .io_inAct(PEs_12_1_io_inAct),
    .io_inWtPS(PEs_12_1_io_inWtPS),
    .io_outWtPS(PEs_12_1_io_outWtPS),
    .io_outAct(PEs_12_1_io_outAct),
    .io_inwtValid(PEs_12_1_io_inwtValid)
  );
  PE PEs_12_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_2_clock),
    .io_inAct(PEs_12_2_io_inAct),
    .io_inWtPS(PEs_12_2_io_inWtPS),
    .io_outWtPS(PEs_12_2_io_outWtPS),
    .io_outAct(PEs_12_2_io_outAct),
    .io_inwtValid(PEs_12_2_io_inwtValid)
  );
  PE PEs_12_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_3_clock),
    .io_inAct(PEs_12_3_io_inAct),
    .io_inWtPS(PEs_12_3_io_inWtPS),
    .io_outWtPS(PEs_12_3_io_outWtPS),
    .io_outAct(PEs_12_3_io_outAct),
    .io_inwtValid(PEs_12_3_io_inwtValid)
  );
  PE PEs_12_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_4_clock),
    .io_inAct(PEs_12_4_io_inAct),
    .io_inWtPS(PEs_12_4_io_inWtPS),
    .io_outWtPS(PEs_12_4_io_outWtPS),
    .io_outAct(PEs_12_4_io_outAct),
    .io_inwtValid(PEs_12_4_io_inwtValid)
  );
  PE PEs_12_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_5_clock),
    .io_inAct(PEs_12_5_io_inAct),
    .io_inWtPS(PEs_12_5_io_inWtPS),
    .io_outWtPS(PEs_12_5_io_outWtPS),
    .io_outAct(PEs_12_5_io_outAct),
    .io_inwtValid(PEs_12_5_io_inwtValid)
  );
  PE PEs_12_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_6_clock),
    .io_inAct(PEs_12_6_io_inAct),
    .io_inWtPS(PEs_12_6_io_inWtPS),
    .io_outWtPS(PEs_12_6_io_outWtPS),
    .io_outAct(PEs_12_6_io_outAct),
    .io_inwtValid(PEs_12_6_io_inwtValid)
  );
  PE PEs_12_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_7_clock),
    .io_inAct(PEs_12_7_io_inAct),
    .io_inWtPS(PEs_12_7_io_inWtPS),
    .io_outWtPS(PEs_12_7_io_outWtPS),
    .io_outAct(PEs_12_7_io_outAct),
    .io_inwtValid(PEs_12_7_io_inwtValid)
  );
  PE PEs_12_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_8_clock),
    .io_inAct(PEs_12_8_io_inAct),
    .io_inWtPS(PEs_12_8_io_inWtPS),
    .io_outWtPS(PEs_12_8_io_outWtPS),
    .io_outAct(PEs_12_8_io_outAct),
    .io_inwtValid(PEs_12_8_io_inwtValid)
  );
  PE PEs_12_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_12_9_clock),
    .io_inAct(PEs_12_9_io_inAct),
    .io_inWtPS(PEs_12_9_io_inWtPS),
    .io_outWtPS(PEs_12_9_io_outWtPS),
    .io_outAct(PEs_12_9_io_outAct),
    .io_inwtValid(PEs_12_9_io_inwtValid)
  );
  PE PEs_13_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_0_clock),
    .io_inAct(PEs_13_0_io_inAct),
    .io_inWtPS(PEs_13_0_io_inWtPS),
    .io_outWtPS(PEs_13_0_io_outWtPS),
    .io_outAct(PEs_13_0_io_outAct),
    .io_inwtValid(PEs_13_0_io_inwtValid)
  );
  PE PEs_13_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_1_clock),
    .io_inAct(PEs_13_1_io_inAct),
    .io_inWtPS(PEs_13_1_io_inWtPS),
    .io_outWtPS(PEs_13_1_io_outWtPS),
    .io_outAct(PEs_13_1_io_outAct),
    .io_inwtValid(PEs_13_1_io_inwtValid)
  );
  PE PEs_13_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_2_clock),
    .io_inAct(PEs_13_2_io_inAct),
    .io_inWtPS(PEs_13_2_io_inWtPS),
    .io_outWtPS(PEs_13_2_io_outWtPS),
    .io_outAct(PEs_13_2_io_outAct),
    .io_inwtValid(PEs_13_2_io_inwtValid)
  );
  PE PEs_13_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_3_clock),
    .io_inAct(PEs_13_3_io_inAct),
    .io_inWtPS(PEs_13_3_io_inWtPS),
    .io_outWtPS(PEs_13_3_io_outWtPS),
    .io_outAct(PEs_13_3_io_outAct),
    .io_inwtValid(PEs_13_3_io_inwtValid)
  );
  PE PEs_13_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_4_clock),
    .io_inAct(PEs_13_4_io_inAct),
    .io_inWtPS(PEs_13_4_io_inWtPS),
    .io_outWtPS(PEs_13_4_io_outWtPS),
    .io_outAct(PEs_13_4_io_outAct),
    .io_inwtValid(PEs_13_4_io_inwtValid)
  );
  PE PEs_13_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_5_clock),
    .io_inAct(PEs_13_5_io_inAct),
    .io_inWtPS(PEs_13_5_io_inWtPS),
    .io_outWtPS(PEs_13_5_io_outWtPS),
    .io_outAct(PEs_13_5_io_outAct),
    .io_inwtValid(PEs_13_5_io_inwtValid)
  );
  PE PEs_13_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_6_clock),
    .io_inAct(PEs_13_6_io_inAct),
    .io_inWtPS(PEs_13_6_io_inWtPS),
    .io_outWtPS(PEs_13_6_io_outWtPS),
    .io_outAct(PEs_13_6_io_outAct),
    .io_inwtValid(PEs_13_6_io_inwtValid)
  );
  PE PEs_13_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_7_clock),
    .io_inAct(PEs_13_7_io_inAct),
    .io_inWtPS(PEs_13_7_io_inWtPS),
    .io_outWtPS(PEs_13_7_io_outWtPS),
    .io_outAct(PEs_13_7_io_outAct),
    .io_inwtValid(PEs_13_7_io_inwtValid)
  );
  PE PEs_13_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_8_clock),
    .io_inAct(PEs_13_8_io_inAct),
    .io_inWtPS(PEs_13_8_io_inWtPS),
    .io_outWtPS(PEs_13_8_io_outWtPS),
    .io_outAct(PEs_13_8_io_outAct),
    .io_inwtValid(PEs_13_8_io_inwtValid)
  );
  PE PEs_13_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_13_9_clock),
    .io_inAct(PEs_13_9_io_inAct),
    .io_inWtPS(PEs_13_9_io_inWtPS),
    .io_outWtPS(PEs_13_9_io_outWtPS),
    .io_outAct(PEs_13_9_io_outAct),
    .io_inwtValid(PEs_13_9_io_inwtValid)
  );
  PE PEs_14_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_0_clock),
    .io_inAct(PEs_14_0_io_inAct),
    .io_inWtPS(PEs_14_0_io_inWtPS),
    .io_outWtPS(PEs_14_0_io_outWtPS),
    .io_outAct(PEs_14_0_io_outAct),
    .io_inwtValid(PEs_14_0_io_inwtValid)
  );
  PE PEs_14_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_1_clock),
    .io_inAct(PEs_14_1_io_inAct),
    .io_inWtPS(PEs_14_1_io_inWtPS),
    .io_outWtPS(PEs_14_1_io_outWtPS),
    .io_outAct(PEs_14_1_io_outAct),
    .io_inwtValid(PEs_14_1_io_inwtValid)
  );
  PE PEs_14_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_2_clock),
    .io_inAct(PEs_14_2_io_inAct),
    .io_inWtPS(PEs_14_2_io_inWtPS),
    .io_outWtPS(PEs_14_2_io_outWtPS),
    .io_outAct(PEs_14_2_io_outAct),
    .io_inwtValid(PEs_14_2_io_inwtValid)
  );
  PE PEs_14_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_3_clock),
    .io_inAct(PEs_14_3_io_inAct),
    .io_inWtPS(PEs_14_3_io_inWtPS),
    .io_outWtPS(PEs_14_3_io_outWtPS),
    .io_outAct(PEs_14_3_io_outAct),
    .io_inwtValid(PEs_14_3_io_inwtValid)
  );
  PE PEs_14_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_4_clock),
    .io_inAct(PEs_14_4_io_inAct),
    .io_inWtPS(PEs_14_4_io_inWtPS),
    .io_outWtPS(PEs_14_4_io_outWtPS),
    .io_outAct(PEs_14_4_io_outAct),
    .io_inwtValid(PEs_14_4_io_inwtValid)
  );
  PE PEs_14_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_5_clock),
    .io_inAct(PEs_14_5_io_inAct),
    .io_inWtPS(PEs_14_5_io_inWtPS),
    .io_outWtPS(PEs_14_5_io_outWtPS),
    .io_outAct(PEs_14_5_io_outAct),
    .io_inwtValid(PEs_14_5_io_inwtValid)
  );
  PE PEs_14_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_6_clock),
    .io_inAct(PEs_14_6_io_inAct),
    .io_inWtPS(PEs_14_6_io_inWtPS),
    .io_outWtPS(PEs_14_6_io_outWtPS),
    .io_outAct(PEs_14_6_io_outAct),
    .io_inwtValid(PEs_14_6_io_inwtValid)
  );
  PE PEs_14_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_7_clock),
    .io_inAct(PEs_14_7_io_inAct),
    .io_inWtPS(PEs_14_7_io_inWtPS),
    .io_outWtPS(PEs_14_7_io_outWtPS),
    .io_outAct(PEs_14_7_io_outAct),
    .io_inwtValid(PEs_14_7_io_inwtValid)
  );
  PE PEs_14_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_8_clock),
    .io_inAct(PEs_14_8_io_inAct),
    .io_inWtPS(PEs_14_8_io_inWtPS),
    .io_outWtPS(PEs_14_8_io_outWtPS),
    .io_outAct(PEs_14_8_io_outAct),
    .io_inwtValid(PEs_14_8_io_inwtValid)
  );
  PE PEs_14_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_14_9_clock),
    .io_inAct(PEs_14_9_io_inAct),
    .io_inWtPS(PEs_14_9_io_inWtPS),
    .io_outWtPS(PEs_14_9_io_outWtPS),
    .io_outAct(PEs_14_9_io_outAct),
    .io_inwtValid(PEs_14_9_io_inwtValid)
  );
  PE PEs_15_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_0_clock),
    .io_inAct(PEs_15_0_io_inAct),
    .io_inWtPS(PEs_15_0_io_inWtPS),
    .io_outWtPS(PEs_15_0_io_outWtPS),
    .io_outAct(PEs_15_0_io_outAct),
    .io_inwtValid(PEs_15_0_io_inwtValid)
  );
  PE PEs_15_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_1_clock),
    .io_inAct(PEs_15_1_io_inAct),
    .io_inWtPS(PEs_15_1_io_inWtPS),
    .io_outWtPS(PEs_15_1_io_outWtPS),
    .io_outAct(PEs_15_1_io_outAct),
    .io_inwtValid(PEs_15_1_io_inwtValid)
  );
  PE PEs_15_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_2_clock),
    .io_inAct(PEs_15_2_io_inAct),
    .io_inWtPS(PEs_15_2_io_inWtPS),
    .io_outWtPS(PEs_15_2_io_outWtPS),
    .io_outAct(PEs_15_2_io_outAct),
    .io_inwtValid(PEs_15_2_io_inwtValid)
  );
  PE PEs_15_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_3_clock),
    .io_inAct(PEs_15_3_io_inAct),
    .io_inWtPS(PEs_15_3_io_inWtPS),
    .io_outWtPS(PEs_15_3_io_outWtPS),
    .io_outAct(PEs_15_3_io_outAct),
    .io_inwtValid(PEs_15_3_io_inwtValid)
  );
  PE PEs_15_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_4_clock),
    .io_inAct(PEs_15_4_io_inAct),
    .io_inWtPS(PEs_15_4_io_inWtPS),
    .io_outWtPS(PEs_15_4_io_outWtPS),
    .io_outAct(PEs_15_4_io_outAct),
    .io_inwtValid(PEs_15_4_io_inwtValid)
  );
  PE PEs_15_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_5_clock),
    .io_inAct(PEs_15_5_io_inAct),
    .io_inWtPS(PEs_15_5_io_inWtPS),
    .io_outWtPS(PEs_15_5_io_outWtPS),
    .io_outAct(PEs_15_5_io_outAct),
    .io_inwtValid(PEs_15_5_io_inwtValid)
  );
  PE PEs_15_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_6_clock),
    .io_inAct(PEs_15_6_io_inAct),
    .io_inWtPS(PEs_15_6_io_inWtPS),
    .io_outWtPS(PEs_15_6_io_outWtPS),
    .io_outAct(PEs_15_6_io_outAct),
    .io_inwtValid(PEs_15_6_io_inwtValid)
  );
  PE PEs_15_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_7_clock),
    .io_inAct(PEs_15_7_io_inAct),
    .io_inWtPS(PEs_15_7_io_inWtPS),
    .io_outWtPS(PEs_15_7_io_outWtPS),
    .io_outAct(PEs_15_7_io_outAct),
    .io_inwtValid(PEs_15_7_io_inwtValid)
  );
  PE PEs_15_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_8_clock),
    .io_inAct(PEs_15_8_io_inAct),
    .io_inWtPS(PEs_15_8_io_inWtPS),
    .io_outWtPS(PEs_15_8_io_outWtPS),
    .io_outAct(PEs_15_8_io_outAct),
    .io_inwtValid(PEs_15_8_io_inwtValid)
  );
  PE PEs_15_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_15_9_clock),
    .io_inAct(PEs_15_9_io_inAct),
    .io_inWtPS(PEs_15_9_io_inWtPS),
    .io_outWtPS(PEs_15_9_io_outWtPS),
    .io_outAct(PEs_15_9_io_outAct),
    .io_inwtValid(PEs_15_9_io_inwtValid)
  );
  PE PEs_16_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_0_clock),
    .io_inAct(PEs_16_0_io_inAct),
    .io_inWtPS(PEs_16_0_io_inWtPS),
    .io_outWtPS(PEs_16_0_io_outWtPS),
    .io_outAct(PEs_16_0_io_outAct),
    .io_inwtValid(PEs_16_0_io_inwtValid)
  );
  PE PEs_16_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_1_clock),
    .io_inAct(PEs_16_1_io_inAct),
    .io_inWtPS(PEs_16_1_io_inWtPS),
    .io_outWtPS(PEs_16_1_io_outWtPS),
    .io_outAct(PEs_16_1_io_outAct),
    .io_inwtValid(PEs_16_1_io_inwtValid)
  );
  PE PEs_16_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_2_clock),
    .io_inAct(PEs_16_2_io_inAct),
    .io_inWtPS(PEs_16_2_io_inWtPS),
    .io_outWtPS(PEs_16_2_io_outWtPS),
    .io_outAct(PEs_16_2_io_outAct),
    .io_inwtValid(PEs_16_2_io_inwtValid)
  );
  PE PEs_16_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_3_clock),
    .io_inAct(PEs_16_3_io_inAct),
    .io_inWtPS(PEs_16_3_io_inWtPS),
    .io_outWtPS(PEs_16_3_io_outWtPS),
    .io_outAct(PEs_16_3_io_outAct),
    .io_inwtValid(PEs_16_3_io_inwtValid)
  );
  PE PEs_16_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_4_clock),
    .io_inAct(PEs_16_4_io_inAct),
    .io_inWtPS(PEs_16_4_io_inWtPS),
    .io_outWtPS(PEs_16_4_io_outWtPS),
    .io_outAct(PEs_16_4_io_outAct),
    .io_inwtValid(PEs_16_4_io_inwtValid)
  );
  PE PEs_16_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_5_clock),
    .io_inAct(PEs_16_5_io_inAct),
    .io_inWtPS(PEs_16_5_io_inWtPS),
    .io_outWtPS(PEs_16_5_io_outWtPS),
    .io_outAct(PEs_16_5_io_outAct),
    .io_inwtValid(PEs_16_5_io_inwtValid)
  );
  PE PEs_16_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_6_clock),
    .io_inAct(PEs_16_6_io_inAct),
    .io_inWtPS(PEs_16_6_io_inWtPS),
    .io_outWtPS(PEs_16_6_io_outWtPS),
    .io_outAct(PEs_16_6_io_outAct),
    .io_inwtValid(PEs_16_6_io_inwtValid)
  );
  PE PEs_16_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_7_clock),
    .io_inAct(PEs_16_7_io_inAct),
    .io_inWtPS(PEs_16_7_io_inWtPS),
    .io_outWtPS(PEs_16_7_io_outWtPS),
    .io_outAct(PEs_16_7_io_outAct),
    .io_inwtValid(PEs_16_7_io_inwtValid)
  );
  PE PEs_16_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_8_clock),
    .io_inAct(PEs_16_8_io_inAct),
    .io_inWtPS(PEs_16_8_io_inWtPS),
    .io_outWtPS(PEs_16_8_io_outWtPS),
    .io_outAct(PEs_16_8_io_outAct),
    .io_inwtValid(PEs_16_8_io_inwtValid)
  );
  PE PEs_16_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_16_9_clock),
    .io_inAct(PEs_16_9_io_inAct),
    .io_inWtPS(PEs_16_9_io_inWtPS),
    .io_outWtPS(PEs_16_9_io_outWtPS),
    .io_outAct(PEs_16_9_io_outAct),
    .io_inwtValid(PEs_16_9_io_inwtValid)
  );
  PE PEs_17_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_0_clock),
    .io_inAct(PEs_17_0_io_inAct),
    .io_inWtPS(PEs_17_0_io_inWtPS),
    .io_outWtPS(PEs_17_0_io_outWtPS),
    .io_outAct(PEs_17_0_io_outAct),
    .io_inwtValid(PEs_17_0_io_inwtValid)
  );
  PE PEs_17_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_1_clock),
    .io_inAct(PEs_17_1_io_inAct),
    .io_inWtPS(PEs_17_1_io_inWtPS),
    .io_outWtPS(PEs_17_1_io_outWtPS),
    .io_outAct(PEs_17_1_io_outAct),
    .io_inwtValid(PEs_17_1_io_inwtValid)
  );
  PE PEs_17_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_2_clock),
    .io_inAct(PEs_17_2_io_inAct),
    .io_inWtPS(PEs_17_2_io_inWtPS),
    .io_outWtPS(PEs_17_2_io_outWtPS),
    .io_outAct(PEs_17_2_io_outAct),
    .io_inwtValid(PEs_17_2_io_inwtValid)
  );
  PE PEs_17_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_3_clock),
    .io_inAct(PEs_17_3_io_inAct),
    .io_inWtPS(PEs_17_3_io_inWtPS),
    .io_outWtPS(PEs_17_3_io_outWtPS),
    .io_outAct(PEs_17_3_io_outAct),
    .io_inwtValid(PEs_17_3_io_inwtValid)
  );
  PE PEs_17_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_4_clock),
    .io_inAct(PEs_17_4_io_inAct),
    .io_inWtPS(PEs_17_4_io_inWtPS),
    .io_outWtPS(PEs_17_4_io_outWtPS),
    .io_outAct(PEs_17_4_io_outAct),
    .io_inwtValid(PEs_17_4_io_inwtValid)
  );
  PE PEs_17_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_5_clock),
    .io_inAct(PEs_17_5_io_inAct),
    .io_inWtPS(PEs_17_5_io_inWtPS),
    .io_outWtPS(PEs_17_5_io_outWtPS),
    .io_outAct(PEs_17_5_io_outAct),
    .io_inwtValid(PEs_17_5_io_inwtValid)
  );
  PE PEs_17_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_6_clock),
    .io_inAct(PEs_17_6_io_inAct),
    .io_inWtPS(PEs_17_6_io_inWtPS),
    .io_outWtPS(PEs_17_6_io_outWtPS),
    .io_outAct(PEs_17_6_io_outAct),
    .io_inwtValid(PEs_17_6_io_inwtValid)
  );
  PE PEs_17_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_7_clock),
    .io_inAct(PEs_17_7_io_inAct),
    .io_inWtPS(PEs_17_7_io_inWtPS),
    .io_outWtPS(PEs_17_7_io_outWtPS),
    .io_outAct(PEs_17_7_io_outAct),
    .io_inwtValid(PEs_17_7_io_inwtValid)
  );
  PE PEs_17_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_8_clock),
    .io_inAct(PEs_17_8_io_inAct),
    .io_inWtPS(PEs_17_8_io_inWtPS),
    .io_outWtPS(PEs_17_8_io_outWtPS),
    .io_outAct(PEs_17_8_io_outAct),
    .io_inwtValid(PEs_17_8_io_inwtValid)
  );
  PE PEs_17_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_17_9_clock),
    .io_inAct(PEs_17_9_io_inAct),
    .io_inWtPS(PEs_17_9_io_inWtPS),
    .io_outWtPS(PEs_17_9_io_outWtPS),
    .io_outAct(PEs_17_9_io_outAct),
    .io_inwtValid(PEs_17_9_io_inwtValid)
  );
  PE PEs_18_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_0_clock),
    .io_inAct(PEs_18_0_io_inAct),
    .io_inWtPS(PEs_18_0_io_inWtPS),
    .io_outWtPS(PEs_18_0_io_outWtPS),
    .io_outAct(PEs_18_0_io_outAct),
    .io_inwtValid(PEs_18_0_io_inwtValid)
  );
  PE PEs_18_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_1_clock),
    .io_inAct(PEs_18_1_io_inAct),
    .io_inWtPS(PEs_18_1_io_inWtPS),
    .io_outWtPS(PEs_18_1_io_outWtPS),
    .io_outAct(PEs_18_1_io_outAct),
    .io_inwtValid(PEs_18_1_io_inwtValid)
  );
  PE PEs_18_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_2_clock),
    .io_inAct(PEs_18_2_io_inAct),
    .io_inWtPS(PEs_18_2_io_inWtPS),
    .io_outWtPS(PEs_18_2_io_outWtPS),
    .io_outAct(PEs_18_2_io_outAct),
    .io_inwtValid(PEs_18_2_io_inwtValid)
  );
  PE PEs_18_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_3_clock),
    .io_inAct(PEs_18_3_io_inAct),
    .io_inWtPS(PEs_18_3_io_inWtPS),
    .io_outWtPS(PEs_18_3_io_outWtPS),
    .io_outAct(PEs_18_3_io_outAct),
    .io_inwtValid(PEs_18_3_io_inwtValid)
  );
  PE PEs_18_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_4_clock),
    .io_inAct(PEs_18_4_io_inAct),
    .io_inWtPS(PEs_18_4_io_inWtPS),
    .io_outWtPS(PEs_18_4_io_outWtPS),
    .io_outAct(PEs_18_4_io_outAct),
    .io_inwtValid(PEs_18_4_io_inwtValid)
  );
  PE PEs_18_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_5_clock),
    .io_inAct(PEs_18_5_io_inAct),
    .io_inWtPS(PEs_18_5_io_inWtPS),
    .io_outWtPS(PEs_18_5_io_outWtPS),
    .io_outAct(PEs_18_5_io_outAct),
    .io_inwtValid(PEs_18_5_io_inwtValid)
  );
  PE PEs_18_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_6_clock),
    .io_inAct(PEs_18_6_io_inAct),
    .io_inWtPS(PEs_18_6_io_inWtPS),
    .io_outWtPS(PEs_18_6_io_outWtPS),
    .io_outAct(PEs_18_6_io_outAct),
    .io_inwtValid(PEs_18_6_io_inwtValid)
  );
  PE PEs_18_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_7_clock),
    .io_inAct(PEs_18_7_io_inAct),
    .io_inWtPS(PEs_18_7_io_inWtPS),
    .io_outWtPS(PEs_18_7_io_outWtPS),
    .io_outAct(PEs_18_7_io_outAct),
    .io_inwtValid(PEs_18_7_io_inwtValid)
  );
  PE PEs_18_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_8_clock),
    .io_inAct(PEs_18_8_io_inAct),
    .io_inWtPS(PEs_18_8_io_inWtPS),
    .io_outWtPS(PEs_18_8_io_outWtPS),
    .io_outAct(PEs_18_8_io_outAct),
    .io_inwtValid(PEs_18_8_io_inwtValid)
  );
  PE PEs_18_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_18_9_clock),
    .io_inAct(PEs_18_9_io_inAct),
    .io_inWtPS(PEs_18_9_io_inWtPS),
    .io_outWtPS(PEs_18_9_io_outWtPS),
    .io_outAct(PEs_18_9_io_outAct),
    .io_inwtValid(PEs_18_9_io_inwtValid)
  );
  PE PEs_19_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_0_clock),
    .io_inAct(PEs_19_0_io_inAct),
    .io_inWtPS(PEs_19_0_io_inWtPS),
    .io_outWtPS(PEs_19_0_io_outWtPS),
    .io_outAct(PEs_19_0_io_outAct),
    .io_inwtValid(PEs_19_0_io_inwtValid)
  );
  PE PEs_19_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_1_clock),
    .io_inAct(PEs_19_1_io_inAct),
    .io_inWtPS(PEs_19_1_io_inWtPS),
    .io_outWtPS(PEs_19_1_io_outWtPS),
    .io_outAct(PEs_19_1_io_outAct),
    .io_inwtValid(PEs_19_1_io_inwtValid)
  );
  PE PEs_19_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_2_clock),
    .io_inAct(PEs_19_2_io_inAct),
    .io_inWtPS(PEs_19_2_io_inWtPS),
    .io_outWtPS(PEs_19_2_io_outWtPS),
    .io_outAct(PEs_19_2_io_outAct),
    .io_inwtValid(PEs_19_2_io_inwtValid)
  );
  PE PEs_19_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_3_clock),
    .io_inAct(PEs_19_3_io_inAct),
    .io_inWtPS(PEs_19_3_io_inWtPS),
    .io_outWtPS(PEs_19_3_io_outWtPS),
    .io_outAct(PEs_19_3_io_outAct),
    .io_inwtValid(PEs_19_3_io_inwtValid)
  );
  PE PEs_19_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_4_clock),
    .io_inAct(PEs_19_4_io_inAct),
    .io_inWtPS(PEs_19_4_io_inWtPS),
    .io_outWtPS(PEs_19_4_io_outWtPS),
    .io_outAct(PEs_19_4_io_outAct),
    .io_inwtValid(PEs_19_4_io_inwtValid)
  );
  PE PEs_19_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_5_clock),
    .io_inAct(PEs_19_5_io_inAct),
    .io_inWtPS(PEs_19_5_io_inWtPS),
    .io_outWtPS(PEs_19_5_io_outWtPS),
    .io_outAct(PEs_19_5_io_outAct),
    .io_inwtValid(PEs_19_5_io_inwtValid)
  );
  PE PEs_19_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_6_clock),
    .io_inAct(PEs_19_6_io_inAct),
    .io_inWtPS(PEs_19_6_io_inWtPS),
    .io_outWtPS(PEs_19_6_io_outWtPS),
    .io_outAct(PEs_19_6_io_outAct),
    .io_inwtValid(PEs_19_6_io_inwtValid)
  );
  PE PEs_19_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_7_clock),
    .io_inAct(PEs_19_7_io_inAct),
    .io_inWtPS(PEs_19_7_io_inWtPS),
    .io_outWtPS(PEs_19_7_io_outWtPS),
    .io_outAct(PEs_19_7_io_outAct),
    .io_inwtValid(PEs_19_7_io_inwtValid)
  );
  PE PEs_19_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_8_clock),
    .io_inAct(PEs_19_8_io_inAct),
    .io_inWtPS(PEs_19_8_io_inWtPS),
    .io_outWtPS(PEs_19_8_io_outWtPS),
    .io_outAct(PEs_19_8_io_outAct),
    .io_inwtValid(PEs_19_8_io_inwtValid)
  );
  PE PEs_19_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_19_9_clock),
    .io_inAct(PEs_19_9_io_inAct),
    .io_inWtPS(PEs_19_9_io_inWtPS),
    .io_outWtPS(PEs_19_9_io_outWtPS),
    .io_outAct(PEs_19_9_io_outAct),
    .io_inwtValid(PEs_19_9_io_inwtValid)
  );
  assign io_outSum_0 = PEs_19_0_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_1 = PEs_19_1_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_2 = PEs_19_2_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_3 = PEs_19_3_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_4 = PEs_19_4_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_5 = PEs_19_5_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_6 = PEs_19_6_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_7 = PEs_19_7_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_8 = PEs_19_8_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_9 = PEs_19_9_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign PEs_0_0_clock = clock;
  assign PEs_0_0_io_inAct = io_inAct_0; // @[SystolicArray.scala 38:44]
  assign PEs_0_0_io_inWtPS = {{24{io_inWeight_0[15]}},io_inWeight_0}; // @[SystolicArray.scala 31:45]
  assign PEs_0_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_1_clock = clock;
  assign PEs_0_1_io_inAct = PEs_0_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_1_io_inWtPS = {{24{io_inWeight_1[15]}},io_inWeight_1}; // @[SystolicArray.scala 31:45]
  assign PEs_0_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_2_clock = clock;
  assign PEs_0_2_io_inAct = PEs_0_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_2_io_inWtPS = {{24{io_inWeight_2[15]}},io_inWeight_2}; // @[SystolicArray.scala 31:45]
  assign PEs_0_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_3_clock = clock;
  assign PEs_0_3_io_inAct = PEs_0_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_3_io_inWtPS = {{24{io_inWeight_3[15]}},io_inWeight_3}; // @[SystolicArray.scala 31:45]
  assign PEs_0_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_4_clock = clock;
  assign PEs_0_4_io_inAct = PEs_0_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_4_io_inWtPS = {{24{io_inWeight_4[15]}},io_inWeight_4}; // @[SystolicArray.scala 31:45]
  assign PEs_0_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_5_clock = clock;
  assign PEs_0_5_io_inAct = PEs_0_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_5_io_inWtPS = {{24{io_inWeight_5[15]}},io_inWeight_5}; // @[SystolicArray.scala 31:45]
  assign PEs_0_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_6_clock = clock;
  assign PEs_0_6_io_inAct = PEs_0_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_6_io_inWtPS = {{24{io_inWeight_6[15]}},io_inWeight_6}; // @[SystolicArray.scala 31:45]
  assign PEs_0_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_7_clock = clock;
  assign PEs_0_7_io_inAct = PEs_0_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_7_io_inWtPS = {{24{io_inWeight_7[15]}},io_inWeight_7}; // @[SystolicArray.scala 31:45]
  assign PEs_0_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_8_clock = clock;
  assign PEs_0_8_io_inAct = PEs_0_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_8_io_inWtPS = {{24{io_inWeight_8[15]}},io_inWeight_8}; // @[SystolicArray.scala 31:45]
  assign PEs_0_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_9_clock = clock;
  assign PEs_0_9_io_inAct = PEs_0_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_9_io_inWtPS = {{24{io_inWeight_9[15]}},io_inWeight_9}; // @[SystolicArray.scala 31:45]
  assign PEs_0_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_0_clock = clock;
  assign PEs_1_0_io_inAct = io_inAct_1; // @[SystolicArray.scala 38:44]
  assign PEs_1_0_io_inWtPS = PEs_0_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_1_clock = clock;
  assign PEs_1_1_io_inAct = PEs_1_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_1_io_inWtPS = PEs_0_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_2_clock = clock;
  assign PEs_1_2_io_inAct = PEs_1_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_2_io_inWtPS = PEs_0_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_3_clock = clock;
  assign PEs_1_3_io_inAct = PEs_1_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_3_io_inWtPS = PEs_0_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_4_clock = clock;
  assign PEs_1_4_io_inAct = PEs_1_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_4_io_inWtPS = PEs_0_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_5_clock = clock;
  assign PEs_1_5_io_inAct = PEs_1_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_5_io_inWtPS = PEs_0_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_6_clock = clock;
  assign PEs_1_6_io_inAct = PEs_1_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_6_io_inWtPS = PEs_0_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_7_clock = clock;
  assign PEs_1_7_io_inAct = PEs_1_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_7_io_inWtPS = PEs_0_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_8_clock = clock;
  assign PEs_1_8_io_inAct = PEs_1_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_8_io_inWtPS = PEs_0_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_9_clock = clock;
  assign PEs_1_9_io_inAct = PEs_1_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_9_io_inWtPS = PEs_0_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_0_clock = clock;
  assign PEs_2_0_io_inAct = io_inAct_2; // @[SystolicArray.scala 38:44]
  assign PEs_2_0_io_inWtPS = PEs_1_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_1_clock = clock;
  assign PEs_2_1_io_inAct = PEs_2_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_1_io_inWtPS = PEs_1_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_2_clock = clock;
  assign PEs_2_2_io_inAct = PEs_2_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_2_io_inWtPS = PEs_1_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_3_clock = clock;
  assign PEs_2_3_io_inAct = PEs_2_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_3_io_inWtPS = PEs_1_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_4_clock = clock;
  assign PEs_2_4_io_inAct = PEs_2_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_4_io_inWtPS = PEs_1_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_5_clock = clock;
  assign PEs_2_5_io_inAct = PEs_2_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_5_io_inWtPS = PEs_1_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_6_clock = clock;
  assign PEs_2_6_io_inAct = PEs_2_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_6_io_inWtPS = PEs_1_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_7_clock = clock;
  assign PEs_2_7_io_inAct = PEs_2_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_7_io_inWtPS = PEs_1_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_8_clock = clock;
  assign PEs_2_8_io_inAct = PEs_2_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_8_io_inWtPS = PEs_1_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_9_clock = clock;
  assign PEs_2_9_io_inAct = PEs_2_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_9_io_inWtPS = PEs_1_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_0_clock = clock;
  assign PEs_3_0_io_inAct = io_inAct_3; // @[SystolicArray.scala 38:44]
  assign PEs_3_0_io_inWtPS = PEs_2_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_1_clock = clock;
  assign PEs_3_1_io_inAct = PEs_3_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_1_io_inWtPS = PEs_2_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_2_clock = clock;
  assign PEs_3_2_io_inAct = PEs_3_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_2_io_inWtPS = PEs_2_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_3_clock = clock;
  assign PEs_3_3_io_inAct = PEs_3_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_3_io_inWtPS = PEs_2_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_4_clock = clock;
  assign PEs_3_4_io_inAct = PEs_3_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_4_io_inWtPS = PEs_2_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_5_clock = clock;
  assign PEs_3_5_io_inAct = PEs_3_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_5_io_inWtPS = PEs_2_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_6_clock = clock;
  assign PEs_3_6_io_inAct = PEs_3_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_6_io_inWtPS = PEs_2_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_7_clock = clock;
  assign PEs_3_7_io_inAct = PEs_3_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_7_io_inWtPS = PEs_2_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_8_clock = clock;
  assign PEs_3_8_io_inAct = PEs_3_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_8_io_inWtPS = PEs_2_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_9_clock = clock;
  assign PEs_3_9_io_inAct = PEs_3_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_9_io_inWtPS = PEs_2_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_0_clock = clock;
  assign PEs_4_0_io_inAct = io_inAct_4; // @[SystolicArray.scala 38:44]
  assign PEs_4_0_io_inWtPS = PEs_3_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_1_clock = clock;
  assign PEs_4_1_io_inAct = PEs_4_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_1_io_inWtPS = PEs_3_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_2_clock = clock;
  assign PEs_4_2_io_inAct = PEs_4_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_2_io_inWtPS = PEs_3_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_3_clock = clock;
  assign PEs_4_3_io_inAct = PEs_4_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_3_io_inWtPS = PEs_3_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_4_clock = clock;
  assign PEs_4_4_io_inAct = PEs_4_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_4_io_inWtPS = PEs_3_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_5_clock = clock;
  assign PEs_4_5_io_inAct = PEs_4_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_5_io_inWtPS = PEs_3_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_6_clock = clock;
  assign PEs_4_6_io_inAct = PEs_4_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_6_io_inWtPS = PEs_3_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_7_clock = clock;
  assign PEs_4_7_io_inAct = PEs_4_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_7_io_inWtPS = PEs_3_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_8_clock = clock;
  assign PEs_4_8_io_inAct = PEs_4_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_8_io_inWtPS = PEs_3_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_9_clock = clock;
  assign PEs_4_9_io_inAct = PEs_4_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_9_io_inWtPS = PEs_3_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_0_clock = clock;
  assign PEs_5_0_io_inAct = io_inAct_5; // @[SystolicArray.scala 38:44]
  assign PEs_5_0_io_inWtPS = PEs_4_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_1_clock = clock;
  assign PEs_5_1_io_inAct = PEs_5_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_1_io_inWtPS = PEs_4_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_2_clock = clock;
  assign PEs_5_2_io_inAct = PEs_5_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_2_io_inWtPS = PEs_4_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_3_clock = clock;
  assign PEs_5_3_io_inAct = PEs_5_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_3_io_inWtPS = PEs_4_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_4_clock = clock;
  assign PEs_5_4_io_inAct = PEs_5_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_4_io_inWtPS = PEs_4_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_5_clock = clock;
  assign PEs_5_5_io_inAct = PEs_5_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_5_io_inWtPS = PEs_4_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_6_clock = clock;
  assign PEs_5_6_io_inAct = PEs_5_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_6_io_inWtPS = PEs_4_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_7_clock = clock;
  assign PEs_5_7_io_inAct = PEs_5_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_7_io_inWtPS = PEs_4_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_8_clock = clock;
  assign PEs_5_8_io_inAct = PEs_5_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_8_io_inWtPS = PEs_4_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_9_clock = clock;
  assign PEs_5_9_io_inAct = PEs_5_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_9_io_inWtPS = PEs_4_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_0_clock = clock;
  assign PEs_6_0_io_inAct = io_inAct_6; // @[SystolicArray.scala 38:44]
  assign PEs_6_0_io_inWtPS = PEs_5_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_1_clock = clock;
  assign PEs_6_1_io_inAct = PEs_6_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_1_io_inWtPS = PEs_5_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_2_clock = clock;
  assign PEs_6_2_io_inAct = PEs_6_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_2_io_inWtPS = PEs_5_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_3_clock = clock;
  assign PEs_6_3_io_inAct = PEs_6_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_3_io_inWtPS = PEs_5_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_4_clock = clock;
  assign PEs_6_4_io_inAct = PEs_6_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_4_io_inWtPS = PEs_5_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_5_clock = clock;
  assign PEs_6_5_io_inAct = PEs_6_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_5_io_inWtPS = PEs_5_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_6_clock = clock;
  assign PEs_6_6_io_inAct = PEs_6_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_6_io_inWtPS = PEs_5_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_7_clock = clock;
  assign PEs_6_7_io_inAct = PEs_6_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_7_io_inWtPS = PEs_5_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_8_clock = clock;
  assign PEs_6_8_io_inAct = PEs_6_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_8_io_inWtPS = PEs_5_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_9_clock = clock;
  assign PEs_6_9_io_inAct = PEs_6_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_9_io_inWtPS = PEs_5_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_0_clock = clock;
  assign PEs_7_0_io_inAct = io_inAct_7; // @[SystolicArray.scala 38:44]
  assign PEs_7_0_io_inWtPS = PEs_6_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_1_clock = clock;
  assign PEs_7_1_io_inAct = PEs_7_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_1_io_inWtPS = PEs_6_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_2_clock = clock;
  assign PEs_7_2_io_inAct = PEs_7_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_2_io_inWtPS = PEs_6_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_3_clock = clock;
  assign PEs_7_3_io_inAct = PEs_7_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_3_io_inWtPS = PEs_6_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_4_clock = clock;
  assign PEs_7_4_io_inAct = PEs_7_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_4_io_inWtPS = PEs_6_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_5_clock = clock;
  assign PEs_7_5_io_inAct = PEs_7_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_5_io_inWtPS = PEs_6_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_6_clock = clock;
  assign PEs_7_6_io_inAct = PEs_7_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_6_io_inWtPS = PEs_6_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_7_clock = clock;
  assign PEs_7_7_io_inAct = PEs_7_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_7_io_inWtPS = PEs_6_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_8_clock = clock;
  assign PEs_7_8_io_inAct = PEs_7_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_8_io_inWtPS = PEs_6_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_9_clock = clock;
  assign PEs_7_9_io_inAct = PEs_7_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_9_io_inWtPS = PEs_6_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_0_clock = clock;
  assign PEs_8_0_io_inAct = io_inAct_8; // @[SystolicArray.scala 38:44]
  assign PEs_8_0_io_inWtPS = PEs_7_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_1_clock = clock;
  assign PEs_8_1_io_inAct = PEs_8_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_1_io_inWtPS = PEs_7_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_2_clock = clock;
  assign PEs_8_2_io_inAct = PEs_8_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_2_io_inWtPS = PEs_7_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_3_clock = clock;
  assign PEs_8_3_io_inAct = PEs_8_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_3_io_inWtPS = PEs_7_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_4_clock = clock;
  assign PEs_8_4_io_inAct = PEs_8_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_4_io_inWtPS = PEs_7_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_5_clock = clock;
  assign PEs_8_5_io_inAct = PEs_8_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_5_io_inWtPS = PEs_7_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_6_clock = clock;
  assign PEs_8_6_io_inAct = PEs_8_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_6_io_inWtPS = PEs_7_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_7_clock = clock;
  assign PEs_8_7_io_inAct = PEs_8_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_7_io_inWtPS = PEs_7_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_8_clock = clock;
  assign PEs_8_8_io_inAct = PEs_8_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_8_io_inWtPS = PEs_7_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_9_clock = clock;
  assign PEs_8_9_io_inAct = PEs_8_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_9_io_inWtPS = PEs_7_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_0_clock = clock;
  assign PEs_9_0_io_inAct = io_inAct_9; // @[SystolicArray.scala 38:44]
  assign PEs_9_0_io_inWtPS = PEs_8_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_1_clock = clock;
  assign PEs_9_1_io_inAct = PEs_9_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_1_io_inWtPS = PEs_8_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_2_clock = clock;
  assign PEs_9_2_io_inAct = PEs_9_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_2_io_inWtPS = PEs_8_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_3_clock = clock;
  assign PEs_9_3_io_inAct = PEs_9_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_3_io_inWtPS = PEs_8_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_4_clock = clock;
  assign PEs_9_4_io_inAct = PEs_9_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_4_io_inWtPS = PEs_8_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_5_clock = clock;
  assign PEs_9_5_io_inAct = PEs_9_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_5_io_inWtPS = PEs_8_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_6_clock = clock;
  assign PEs_9_6_io_inAct = PEs_9_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_6_io_inWtPS = PEs_8_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_7_clock = clock;
  assign PEs_9_7_io_inAct = PEs_9_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_7_io_inWtPS = PEs_8_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_8_clock = clock;
  assign PEs_9_8_io_inAct = PEs_9_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_8_io_inWtPS = PEs_8_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_9_clock = clock;
  assign PEs_9_9_io_inAct = PEs_9_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_9_io_inWtPS = PEs_8_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_0_clock = clock;
  assign PEs_10_0_io_inAct = io_inAct_10; // @[SystolicArray.scala 38:44]
  assign PEs_10_0_io_inWtPS = PEs_9_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_1_clock = clock;
  assign PEs_10_1_io_inAct = PEs_10_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_1_io_inWtPS = PEs_9_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_2_clock = clock;
  assign PEs_10_2_io_inAct = PEs_10_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_2_io_inWtPS = PEs_9_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_3_clock = clock;
  assign PEs_10_3_io_inAct = PEs_10_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_3_io_inWtPS = PEs_9_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_4_clock = clock;
  assign PEs_10_4_io_inAct = PEs_10_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_4_io_inWtPS = PEs_9_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_5_clock = clock;
  assign PEs_10_5_io_inAct = PEs_10_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_5_io_inWtPS = PEs_9_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_6_clock = clock;
  assign PEs_10_6_io_inAct = PEs_10_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_6_io_inWtPS = PEs_9_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_7_clock = clock;
  assign PEs_10_7_io_inAct = PEs_10_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_7_io_inWtPS = PEs_9_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_8_clock = clock;
  assign PEs_10_8_io_inAct = PEs_10_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_8_io_inWtPS = PEs_9_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_10_9_clock = clock;
  assign PEs_10_9_io_inAct = PEs_10_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_10_9_io_inWtPS = PEs_9_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_10_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_0_clock = clock;
  assign PEs_11_0_io_inAct = io_inAct_11; // @[SystolicArray.scala 38:44]
  assign PEs_11_0_io_inWtPS = PEs_10_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_1_clock = clock;
  assign PEs_11_1_io_inAct = PEs_11_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_1_io_inWtPS = PEs_10_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_2_clock = clock;
  assign PEs_11_2_io_inAct = PEs_11_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_2_io_inWtPS = PEs_10_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_3_clock = clock;
  assign PEs_11_3_io_inAct = PEs_11_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_3_io_inWtPS = PEs_10_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_4_clock = clock;
  assign PEs_11_4_io_inAct = PEs_11_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_4_io_inWtPS = PEs_10_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_5_clock = clock;
  assign PEs_11_5_io_inAct = PEs_11_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_5_io_inWtPS = PEs_10_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_6_clock = clock;
  assign PEs_11_6_io_inAct = PEs_11_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_6_io_inWtPS = PEs_10_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_7_clock = clock;
  assign PEs_11_7_io_inAct = PEs_11_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_7_io_inWtPS = PEs_10_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_8_clock = clock;
  assign PEs_11_8_io_inAct = PEs_11_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_8_io_inWtPS = PEs_10_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_11_9_clock = clock;
  assign PEs_11_9_io_inAct = PEs_11_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_11_9_io_inWtPS = PEs_10_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_11_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_0_clock = clock;
  assign PEs_12_0_io_inAct = io_inAct_12; // @[SystolicArray.scala 38:44]
  assign PEs_12_0_io_inWtPS = PEs_11_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_1_clock = clock;
  assign PEs_12_1_io_inAct = PEs_12_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_1_io_inWtPS = PEs_11_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_2_clock = clock;
  assign PEs_12_2_io_inAct = PEs_12_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_2_io_inWtPS = PEs_11_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_3_clock = clock;
  assign PEs_12_3_io_inAct = PEs_12_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_3_io_inWtPS = PEs_11_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_4_clock = clock;
  assign PEs_12_4_io_inAct = PEs_12_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_4_io_inWtPS = PEs_11_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_5_clock = clock;
  assign PEs_12_5_io_inAct = PEs_12_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_5_io_inWtPS = PEs_11_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_6_clock = clock;
  assign PEs_12_6_io_inAct = PEs_12_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_6_io_inWtPS = PEs_11_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_7_clock = clock;
  assign PEs_12_7_io_inAct = PEs_12_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_7_io_inWtPS = PEs_11_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_8_clock = clock;
  assign PEs_12_8_io_inAct = PEs_12_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_8_io_inWtPS = PEs_11_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_12_9_clock = clock;
  assign PEs_12_9_io_inAct = PEs_12_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_12_9_io_inWtPS = PEs_11_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_12_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_0_clock = clock;
  assign PEs_13_0_io_inAct = io_inAct_13; // @[SystolicArray.scala 38:44]
  assign PEs_13_0_io_inWtPS = PEs_12_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_1_clock = clock;
  assign PEs_13_1_io_inAct = PEs_13_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_1_io_inWtPS = PEs_12_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_2_clock = clock;
  assign PEs_13_2_io_inAct = PEs_13_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_2_io_inWtPS = PEs_12_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_3_clock = clock;
  assign PEs_13_3_io_inAct = PEs_13_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_3_io_inWtPS = PEs_12_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_4_clock = clock;
  assign PEs_13_4_io_inAct = PEs_13_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_4_io_inWtPS = PEs_12_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_5_clock = clock;
  assign PEs_13_5_io_inAct = PEs_13_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_5_io_inWtPS = PEs_12_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_6_clock = clock;
  assign PEs_13_6_io_inAct = PEs_13_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_6_io_inWtPS = PEs_12_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_7_clock = clock;
  assign PEs_13_7_io_inAct = PEs_13_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_7_io_inWtPS = PEs_12_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_8_clock = clock;
  assign PEs_13_8_io_inAct = PEs_13_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_8_io_inWtPS = PEs_12_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_13_9_clock = clock;
  assign PEs_13_9_io_inAct = PEs_13_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_13_9_io_inWtPS = PEs_12_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_13_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_0_clock = clock;
  assign PEs_14_0_io_inAct = io_inAct_14; // @[SystolicArray.scala 38:44]
  assign PEs_14_0_io_inWtPS = PEs_13_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_1_clock = clock;
  assign PEs_14_1_io_inAct = PEs_14_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_1_io_inWtPS = PEs_13_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_2_clock = clock;
  assign PEs_14_2_io_inAct = PEs_14_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_2_io_inWtPS = PEs_13_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_3_clock = clock;
  assign PEs_14_3_io_inAct = PEs_14_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_3_io_inWtPS = PEs_13_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_4_clock = clock;
  assign PEs_14_4_io_inAct = PEs_14_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_4_io_inWtPS = PEs_13_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_5_clock = clock;
  assign PEs_14_5_io_inAct = PEs_14_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_5_io_inWtPS = PEs_13_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_6_clock = clock;
  assign PEs_14_6_io_inAct = PEs_14_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_6_io_inWtPS = PEs_13_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_7_clock = clock;
  assign PEs_14_7_io_inAct = PEs_14_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_7_io_inWtPS = PEs_13_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_8_clock = clock;
  assign PEs_14_8_io_inAct = PEs_14_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_8_io_inWtPS = PEs_13_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_14_9_clock = clock;
  assign PEs_14_9_io_inAct = PEs_14_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_14_9_io_inWtPS = PEs_13_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_14_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_0_clock = clock;
  assign PEs_15_0_io_inAct = io_inAct_15; // @[SystolicArray.scala 38:44]
  assign PEs_15_0_io_inWtPS = PEs_14_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_1_clock = clock;
  assign PEs_15_1_io_inAct = PEs_15_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_1_io_inWtPS = PEs_14_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_2_clock = clock;
  assign PEs_15_2_io_inAct = PEs_15_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_2_io_inWtPS = PEs_14_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_3_clock = clock;
  assign PEs_15_3_io_inAct = PEs_15_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_3_io_inWtPS = PEs_14_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_4_clock = clock;
  assign PEs_15_4_io_inAct = PEs_15_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_4_io_inWtPS = PEs_14_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_5_clock = clock;
  assign PEs_15_5_io_inAct = PEs_15_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_5_io_inWtPS = PEs_14_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_6_clock = clock;
  assign PEs_15_6_io_inAct = PEs_15_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_6_io_inWtPS = PEs_14_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_7_clock = clock;
  assign PEs_15_7_io_inAct = PEs_15_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_7_io_inWtPS = PEs_14_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_8_clock = clock;
  assign PEs_15_8_io_inAct = PEs_15_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_8_io_inWtPS = PEs_14_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_15_9_clock = clock;
  assign PEs_15_9_io_inAct = PEs_15_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_15_9_io_inWtPS = PEs_14_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_15_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_0_clock = clock;
  assign PEs_16_0_io_inAct = io_inAct_16; // @[SystolicArray.scala 38:44]
  assign PEs_16_0_io_inWtPS = PEs_15_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_1_clock = clock;
  assign PEs_16_1_io_inAct = PEs_16_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_1_io_inWtPS = PEs_15_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_2_clock = clock;
  assign PEs_16_2_io_inAct = PEs_16_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_2_io_inWtPS = PEs_15_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_3_clock = clock;
  assign PEs_16_3_io_inAct = PEs_16_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_3_io_inWtPS = PEs_15_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_4_clock = clock;
  assign PEs_16_4_io_inAct = PEs_16_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_4_io_inWtPS = PEs_15_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_5_clock = clock;
  assign PEs_16_5_io_inAct = PEs_16_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_5_io_inWtPS = PEs_15_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_6_clock = clock;
  assign PEs_16_6_io_inAct = PEs_16_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_6_io_inWtPS = PEs_15_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_7_clock = clock;
  assign PEs_16_7_io_inAct = PEs_16_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_7_io_inWtPS = PEs_15_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_8_clock = clock;
  assign PEs_16_8_io_inAct = PEs_16_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_8_io_inWtPS = PEs_15_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_16_9_clock = clock;
  assign PEs_16_9_io_inAct = PEs_16_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_16_9_io_inWtPS = PEs_15_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_16_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_0_clock = clock;
  assign PEs_17_0_io_inAct = io_inAct_17; // @[SystolicArray.scala 38:44]
  assign PEs_17_0_io_inWtPS = PEs_16_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_1_clock = clock;
  assign PEs_17_1_io_inAct = PEs_17_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_1_io_inWtPS = PEs_16_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_2_clock = clock;
  assign PEs_17_2_io_inAct = PEs_17_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_2_io_inWtPS = PEs_16_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_3_clock = clock;
  assign PEs_17_3_io_inAct = PEs_17_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_3_io_inWtPS = PEs_16_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_4_clock = clock;
  assign PEs_17_4_io_inAct = PEs_17_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_4_io_inWtPS = PEs_16_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_5_clock = clock;
  assign PEs_17_5_io_inAct = PEs_17_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_5_io_inWtPS = PEs_16_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_6_clock = clock;
  assign PEs_17_6_io_inAct = PEs_17_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_6_io_inWtPS = PEs_16_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_7_clock = clock;
  assign PEs_17_7_io_inAct = PEs_17_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_7_io_inWtPS = PEs_16_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_8_clock = clock;
  assign PEs_17_8_io_inAct = PEs_17_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_8_io_inWtPS = PEs_16_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_17_9_clock = clock;
  assign PEs_17_9_io_inAct = PEs_17_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_17_9_io_inWtPS = PEs_16_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_17_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_0_clock = clock;
  assign PEs_18_0_io_inAct = io_inAct_18; // @[SystolicArray.scala 38:44]
  assign PEs_18_0_io_inWtPS = PEs_17_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_1_clock = clock;
  assign PEs_18_1_io_inAct = PEs_18_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_1_io_inWtPS = PEs_17_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_2_clock = clock;
  assign PEs_18_2_io_inAct = PEs_18_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_2_io_inWtPS = PEs_17_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_3_clock = clock;
  assign PEs_18_3_io_inAct = PEs_18_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_3_io_inWtPS = PEs_17_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_4_clock = clock;
  assign PEs_18_4_io_inAct = PEs_18_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_4_io_inWtPS = PEs_17_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_5_clock = clock;
  assign PEs_18_5_io_inAct = PEs_18_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_5_io_inWtPS = PEs_17_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_6_clock = clock;
  assign PEs_18_6_io_inAct = PEs_18_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_6_io_inWtPS = PEs_17_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_7_clock = clock;
  assign PEs_18_7_io_inAct = PEs_18_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_7_io_inWtPS = PEs_17_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_8_clock = clock;
  assign PEs_18_8_io_inAct = PEs_18_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_8_io_inWtPS = PEs_17_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_18_9_clock = clock;
  assign PEs_18_9_io_inAct = PEs_18_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_18_9_io_inWtPS = PEs_17_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_18_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_0_clock = clock;
  assign PEs_19_0_io_inAct = io_inAct_19; // @[SystolicArray.scala 38:44]
  assign PEs_19_0_io_inWtPS = PEs_18_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_1_clock = clock;
  assign PEs_19_1_io_inAct = PEs_19_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_1_io_inWtPS = PEs_18_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_2_clock = clock;
  assign PEs_19_2_io_inAct = PEs_19_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_2_io_inWtPS = PEs_18_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_3_clock = clock;
  assign PEs_19_3_io_inAct = PEs_19_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_3_io_inWtPS = PEs_18_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_4_clock = clock;
  assign PEs_19_4_io_inAct = PEs_19_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_4_io_inWtPS = PEs_18_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_5_clock = clock;
  assign PEs_19_5_io_inAct = PEs_19_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_5_io_inWtPS = PEs_18_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_6_clock = clock;
  assign PEs_19_6_io_inAct = PEs_19_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_6_io_inWtPS = PEs_18_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_7_clock = clock;
  assign PEs_19_7_io_inAct = PEs_19_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_7_io_inWtPS = PEs_18_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_8_clock = clock;
  assign PEs_19_8_io_inAct = PEs_19_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_8_io_inWtPS = PEs_18_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_19_9_clock = clock;
  assign PEs_19_9_io_inAct = PEs_19_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_19_9_io_inWtPS = PEs_18_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_19_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  always @(posedge clock) begin
    validReg <= io_inwtValid; // @[SystolicArray.scala 22:25]
  end
endmodule
module SystolicArray_1(
  input         clock,
  input  [15:0] io_inAct_0,
  input  [15:0] io_inAct_1,
  input  [15:0] io_inAct_2,
  input  [15:0] io_inAct_3,
  input  [15:0] io_inAct_4,
  input  [15:0] io_inAct_5,
  input  [15:0] io_inAct_6,
  input  [15:0] io_inAct_7,
  input  [15:0] io_inAct_8,
  input  [15:0] io_inAct_9,
  input  [15:0] io_inWeight_0,
  input  [15:0] io_inWeight_1,
  input  [15:0] io_inWeight_2,
  input  [15:0] io_inWeight_3,
  input  [15:0] io_inWeight_4,
  input  [15:0] io_inWeight_5,
  input  [15:0] io_inWeight_6,
  input  [15:0] io_inWeight_7,
  input  [15:0] io_inWeight_8,
  input  [15:0] io_inWeight_9,
  output [39:0] io_outSum_0,
  output [39:0] io_outSum_1,
  output [39:0] io_outSum_2,
  output [39:0] io_outSum_3,
  output [39:0] io_outSum_4,
  output [39:0] io_outSum_5,
  output [39:0] io_outSum_6,
  output [39:0] io_outSum_7,
  output [39:0] io_outSum_8,
  output [39:0] io_outSum_9,
  input         io_inwtValid
);
  wire  PEs_0_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_8_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_8_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_8_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_8_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_8_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_8_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_9_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_9_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_9_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_9_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_9_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_9_io_inwtValid; // @[SystolicArray.scala 18:65]
  reg  validReg; // @[SystolicArray.scala 22:25]
  PE PEs_0_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_0_clock),
    .io_inAct(PEs_0_0_io_inAct),
    .io_inWtPS(PEs_0_0_io_inWtPS),
    .io_outWtPS(PEs_0_0_io_outWtPS),
    .io_outAct(PEs_0_0_io_outAct),
    .io_inwtValid(PEs_0_0_io_inwtValid)
  );
  PE PEs_0_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_1_clock),
    .io_inAct(PEs_0_1_io_inAct),
    .io_inWtPS(PEs_0_1_io_inWtPS),
    .io_outWtPS(PEs_0_1_io_outWtPS),
    .io_outAct(PEs_0_1_io_outAct),
    .io_inwtValid(PEs_0_1_io_inwtValid)
  );
  PE PEs_0_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_2_clock),
    .io_inAct(PEs_0_2_io_inAct),
    .io_inWtPS(PEs_0_2_io_inWtPS),
    .io_outWtPS(PEs_0_2_io_outWtPS),
    .io_outAct(PEs_0_2_io_outAct),
    .io_inwtValid(PEs_0_2_io_inwtValid)
  );
  PE PEs_0_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_3_clock),
    .io_inAct(PEs_0_3_io_inAct),
    .io_inWtPS(PEs_0_3_io_inWtPS),
    .io_outWtPS(PEs_0_3_io_outWtPS),
    .io_outAct(PEs_0_3_io_outAct),
    .io_inwtValid(PEs_0_3_io_inwtValid)
  );
  PE PEs_0_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_4_clock),
    .io_inAct(PEs_0_4_io_inAct),
    .io_inWtPS(PEs_0_4_io_inWtPS),
    .io_outWtPS(PEs_0_4_io_outWtPS),
    .io_outAct(PEs_0_4_io_outAct),
    .io_inwtValid(PEs_0_4_io_inwtValid)
  );
  PE PEs_0_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_5_clock),
    .io_inAct(PEs_0_5_io_inAct),
    .io_inWtPS(PEs_0_5_io_inWtPS),
    .io_outWtPS(PEs_0_5_io_outWtPS),
    .io_outAct(PEs_0_5_io_outAct),
    .io_inwtValid(PEs_0_5_io_inwtValid)
  );
  PE PEs_0_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_6_clock),
    .io_inAct(PEs_0_6_io_inAct),
    .io_inWtPS(PEs_0_6_io_inWtPS),
    .io_outWtPS(PEs_0_6_io_outWtPS),
    .io_outAct(PEs_0_6_io_outAct),
    .io_inwtValid(PEs_0_6_io_inwtValid)
  );
  PE PEs_0_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_7_clock),
    .io_inAct(PEs_0_7_io_inAct),
    .io_inWtPS(PEs_0_7_io_inWtPS),
    .io_outWtPS(PEs_0_7_io_outWtPS),
    .io_outAct(PEs_0_7_io_outAct),
    .io_inwtValid(PEs_0_7_io_inwtValid)
  );
  PE PEs_0_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_8_clock),
    .io_inAct(PEs_0_8_io_inAct),
    .io_inWtPS(PEs_0_8_io_inWtPS),
    .io_outWtPS(PEs_0_8_io_outWtPS),
    .io_outAct(PEs_0_8_io_outAct),
    .io_inwtValid(PEs_0_8_io_inwtValid)
  );
  PE PEs_0_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_9_clock),
    .io_inAct(PEs_0_9_io_inAct),
    .io_inWtPS(PEs_0_9_io_inWtPS),
    .io_outWtPS(PEs_0_9_io_outWtPS),
    .io_outAct(PEs_0_9_io_outAct),
    .io_inwtValid(PEs_0_9_io_inwtValid)
  );
  PE PEs_1_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_0_clock),
    .io_inAct(PEs_1_0_io_inAct),
    .io_inWtPS(PEs_1_0_io_inWtPS),
    .io_outWtPS(PEs_1_0_io_outWtPS),
    .io_outAct(PEs_1_0_io_outAct),
    .io_inwtValid(PEs_1_0_io_inwtValid)
  );
  PE PEs_1_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_1_clock),
    .io_inAct(PEs_1_1_io_inAct),
    .io_inWtPS(PEs_1_1_io_inWtPS),
    .io_outWtPS(PEs_1_1_io_outWtPS),
    .io_outAct(PEs_1_1_io_outAct),
    .io_inwtValid(PEs_1_1_io_inwtValid)
  );
  PE PEs_1_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_2_clock),
    .io_inAct(PEs_1_2_io_inAct),
    .io_inWtPS(PEs_1_2_io_inWtPS),
    .io_outWtPS(PEs_1_2_io_outWtPS),
    .io_outAct(PEs_1_2_io_outAct),
    .io_inwtValid(PEs_1_2_io_inwtValid)
  );
  PE PEs_1_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_3_clock),
    .io_inAct(PEs_1_3_io_inAct),
    .io_inWtPS(PEs_1_3_io_inWtPS),
    .io_outWtPS(PEs_1_3_io_outWtPS),
    .io_outAct(PEs_1_3_io_outAct),
    .io_inwtValid(PEs_1_3_io_inwtValid)
  );
  PE PEs_1_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_4_clock),
    .io_inAct(PEs_1_4_io_inAct),
    .io_inWtPS(PEs_1_4_io_inWtPS),
    .io_outWtPS(PEs_1_4_io_outWtPS),
    .io_outAct(PEs_1_4_io_outAct),
    .io_inwtValid(PEs_1_4_io_inwtValid)
  );
  PE PEs_1_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_5_clock),
    .io_inAct(PEs_1_5_io_inAct),
    .io_inWtPS(PEs_1_5_io_inWtPS),
    .io_outWtPS(PEs_1_5_io_outWtPS),
    .io_outAct(PEs_1_5_io_outAct),
    .io_inwtValid(PEs_1_5_io_inwtValid)
  );
  PE PEs_1_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_6_clock),
    .io_inAct(PEs_1_6_io_inAct),
    .io_inWtPS(PEs_1_6_io_inWtPS),
    .io_outWtPS(PEs_1_6_io_outWtPS),
    .io_outAct(PEs_1_6_io_outAct),
    .io_inwtValid(PEs_1_6_io_inwtValid)
  );
  PE PEs_1_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_7_clock),
    .io_inAct(PEs_1_7_io_inAct),
    .io_inWtPS(PEs_1_7_io_inWtPS),
    .io_outWtPS(PEs_1_7_io_outWtPS),
    .io_outAct(PEs_1_7_io_outAct),
    .io_inwtValid(PEs_1_7_io_inwtValid)
  );
  PE PEs_1_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_8_clock),
    .io_inAct(PEs_1_8_io_inAct),
    .io_inWtPS(PEs_1_8_io_inWtPS),
    .io_outWtPS(PEs_1_8_io_outWtPS),
    .io_outAct(PEs_1_8_io_outAct),
    .io_inwtValid(PEs_1_8_io_inwtValid)
  );
  PE PEs_1_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_9_clock),
    .io_inAct(PEs_1_9_io_inAct),
    .io_inWtPS(PEs_1_9_io_inWtPS),
    .io_outWtPS(PEs_1_9_io_outWtPS),
    .io_outAct(PEs_1_9_io_outAct),
    .io_inwtValid(PEs_1_9_io_inwtValid)
  );
  PE PEs_2_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_0_clock),
    .io_inAct(PEs_2_0_io_inAct),
    .io_inWtPS(PEs_2_0_io_inWtPS),
    .io_outWtPS(PEs_2_0_io_outWtPS),
    .io_outAct(PEs_2_0_io_outAct),
    .io_inwtValid(PEs_2_0_io_inwtValid)
  );
  PE PEs_2_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_1_clock),
    .io_inAct(PEs_2_1_io_inAct),
    .io_inWtPS(PEs_2_1_io_inWtPS),
    .io_outWtPS(PEs_2_1_io_outWtPS),
    .io_outAct(PEs_2_1_io_outAct),
    .io_inwtValid(PEs_2_1_io_inwtValid)
  );
  PE PEs_2_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_2_clock),
    .io_inAct(PEs_2_2_io_inAct),
    .io_inWtPS(PEs_2_2_io_inWtPS),
    .io_outWtPS(PEs_2_2_io_outWtPS),
    .io_outAct(PEs_2_2_io_outAct),
    .io_inwtValid(PEs_2_2_io_inwtValid)
  );
  PE PEs_2_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_3_clock),
    .io_inAct(PEs_2_3_io_inAct),
    .io_inWtPS(PEs_2_3_io_inWtPS),
    .io_outWtPS(PEs_2_3_io_outWtPS),
    .io_outAct(PEs_2_3_io_outAct),
    .io_inwtValid(PEs_2_3_io_inwtValid)
  );
  PE PEs_2_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_4_clock),
    .io_inAct(PEs_2_4_io_inAct),
    .io_inWtPS(PEs_2_4_io_inWtPS),
    .io_outWtPS(PEs_2_4_io_outWtPS),
    .io_outAct(PEs_2_4_io_outAct),
    .io_inwtValid(PEs_2_4_io_inwtValid)
  );
  PE PEs_2_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_5_clock),
    .io_inAct(PEs_2_5_io_inAct),
    .io_inWtPS(PEs_2_5_io_inWtPS),
    .io_outWtPS(PEs_2_5_io_outWtPS),
    .io_outAct(PEs_2_5_io_outAct),
    .io_inwtValid(PEs_2_5_io_inwtValid)
  );
  PE PEs_2_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_6_clock),
    .io_inAct(PEs_2_6_io_inAct),
    .io_inWtPS(PEs_2_6_io_inWtPS),
    .io_outWtPS(PEs_2_6_io_outWtPS),
    .io_outAct(PEs_2_6_io_outAct),
    .io_inwtValid(PEs_2_6_io_inwtValid)
  );
  PE PEs_2_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_7_clock),
    .io_inAct(PEs_2_7_io_inAct),
    .io_inWtPS(PEs_2_7_io_inWtPS),
    .io_outWtPS(PEs_2_7_io_outWtPS),
    .io_outAct(PEs_2_7_io_outAct),
    .io_inwtValid(PEs_2_7_io_inwtValid)
  );
  PE PEs_2_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_8_clock),
    .io_inAct(PEs_2_8_io_inAct),
    .io_inWtPS(PEs_2_8_io_inWtPS),
    .io_outWtPS(PEs_2_8_io_outWtPS),
    .io_outAct(PEs_2_8_io_outAct),
    .io_inwtValid(PEs_2_8_io_inwtValid)
  );
  PE PEs_2_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_9_clock),
    .io_inAct(PEs_2_9_io_inAct),
    .io_inWtPS(PEs_2_9_io_inWtPS),
    .io_outWtPS(PEs_2_9_io_outWtPS),
    .io_outAct(PEs_2_9_io_outAct),
    .io_inwtValid(PEs_2_9_io_inwtValid)
  );
  PE PEs_3_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_0_clock),
    .io_inAct(PEs_3_0_io_inAct),
    .io_inWtPS(PEs_3_0_io_inWtPS),
    .io_outWtPS(PEs_3_0_io_outWtPS),
    .io_outAct(PEs_3_0_io_outAct),
    .io_inwtValid(PEs_3_0_io_inwtValid)
  );
  PE PEs_3_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_1_clock),
    .io_inAct(PEs_3_1_io_inAct),
    .io_inWtPS(PEs_3_1_io_inWtPS),
    .io_outWtPS(PEs_3_1_io_outWtPS),
    .io_outAct(PEs_3_1_io_outAct),
    .io_inwtValid(PEs_3_1_io_inwtValid)
  );
  PE PEs_3_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_2_clock),
    .io_inAct(PEs_3_2_io_inAct),
    .io_inWtPS(PEs_3_2_io_inWtPS),
    .io_outWtPS(PEs_3_2_io_outWtPS),
    .io_outAct(PEs_3_2_io_outAct),
    .io_inwtValid(PEs_3_2_io_inwtValid)
  );
  PE PEs_3_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_3_clock),
    .io_inAct(PEs_3_3_io_inAct),
    .io_inWtPS(PEs_3_3_io_inWtPS),
    .io_outWtPS(PEs_3_3_io_outWtPS),
    .io_outAct(PEs_3_3_io_outAct),
    .io_inwtValid(PEs_3_3_io_inwtValid)
  );
  PE PEs_3_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_4_clock),
    .io_inAct(PEs_3_4_io_inAct),
    .io_inWtPS(PEs_3_4_io_inWtPS),
    .io_outWtPS(PEs_3_4_io_outWtPS),
    .io_outAct(PEs_3_4_io_outAct),
    .io_inwtValid(PEs_3_4_io_inwtValid)
  );
  PE PEs_3_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_5_clock),
    .io_inAct(PEs_3_5_io_inAct),
    .io_inWtPS(PEs_3_5_io_inWtPS),
    .io_outWtPS(PEs_3_5_io_outWtPS),
    .io_outAct(PEs_3_5_io_outAct),
    .io_inwtValid(PEs_3_5_io_inwtValid)
  );
  PE PEs_3_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_6_clock),
    .io_inAct(PEs_3_6_io_inAct),
    .io_inWtPS(PEs_3_6_io_inWtPS),
    .io_outWtPS(PEs_3_6_io_outWtPS),
    .io_outAct(PEs_3_6_io_outAct),
    .io_inwtValid(PEs_3_6_io_inwtValid)
  );
  PE PEs_3_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_7_clock),
    .io_inAct(PEs_3_7_io_inAct),
    .io_inWtPS(PEs_3_7_io_inWtPS),
    .io_outWtPS(PEs_3_7_io_outWtPS),
    .io_outAct(PEs_3_7_io_outAct),
    .io_inwtValid(PEs_3_7_io_inwtValid)
  );
  PE PEs_3_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_8_clock),
    .io_inAct(PEs_3_8_io_inAct),
    .io_inWtPS(PEs_3_8_io_inWtPS),
    .io_outWtPS(PEs_3_8_io_outWtPS),
    .io_outAct(PEs_3_8_io_outAct),
    .io_inwtValid(PEs_3_8_io_inwtValid)
  );
  PE PEs_3_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_9_clock),
    .io_inAct(PEs_3_9_io_inAct),
    .io_inWtPS(PEs_3_9_io_inWtPS),
    .io_outWtPS(PEs_3_9_io_outWtPS),
    .io_outAct(PEs_3_9_io_outAct),
    .io_inwtValid(PEs_3_9_io_inwtValid)
  );
  PE PEs_4_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_0_clock),
    .io_inAct(PEs_4_0_io_inAct),
    .io_inWtPS(PEs_4_0_io_inWtPS),
    .io_outWtPS(PEs_4_0_io_outWtPS),
    .io_outAct(PEs_4_0_io_outAct),
    .io_inwtValid(PEs_4_0_io_inwtValid)
  );
  PE PEs_4_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_1_clock),
    .io_inAct(PEs_4_1_io_inAct),
    .io_inWtPS(PEs_4_1_io_inWtPS),
    .io_outWtPS(PEs_4_1_io_outWtPS),
    .io_outAct(PEs_4_1_io_outAct),
    .io_inwtValid(PEs_4_1_io_inwtValid)
  );
  PE PEs_4_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_2_clock),
    .io_inAct(PEs_4_2_io_inAct),
    .io_inWtPS(PEs_4_2_io_inWtPS),
    .io_outWtPS(PEs_4_2_io_outWtPS),
    .io_outAct(PEs_4_2_io_outAct),
    .io_inwtValid(PEs_4_2_io_inwtValid)
  );
  PE PEs_4_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_3_clock),
    .io_inAct(PEs_4_3_io_inAct),
    .io_inWtPS(PEs_4_3_io_inWtPS),
    .io_outWtPS(PEs_4_3_io_outWtPS),
    .io_outAct(PEs_4_3_io_outAct),
    .io_inwtValid(PEs_4_3_io_inwtValid)
  );
  PE PEs_4_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_4_clock),
    .io_inAct(PEs_4_4_io_inAct),
    .io_inWtPS(PEs_4_4_io_inWtPS),
    .io_outWtPS(PEs_4_4_io_outWtPS),
    .io_outAct(PEs_4_4_io_outAct),
    .io_inwtValid(PEs_4_4_io_inwtValid)
  );
  PE PEs_4_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_5_clock),
    .io_inAct(PEs_4_5_io_inAct),
    .io_inWtPS(PEs_4_5_io_inWtPS),
    .io_outWtPS(PEs_4_5_io_outWtPS),
    .io_outAct(PEs_4_5_io_outAct),
    .io_inwtValid(PEs_4_5_io_inwtValid)
  );
  PE PEs_4_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_6_clock),
    .io_inAct(PEs_4_6_io_inAct),
    .io_inWtPS(PEs_4_6_io_inWtPS),
    .io_outWtPS(PEs_4_6_io_outWtPS),
    .io_outAct(PEs_4_6_io_outAct),
    .io_inwtValid(PEs_4_6_io_inwtValid)
  );
  PE PEs_4_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_7_clock),
    .io_inAct(PEs_4_7_io_inAct),
    .io_inWtPS(PEs_4_7_io_inWtPS),
    .io_outWtPS(PEs_4_7_io_outWtPS),
    .io_outAct(PEs_4_7_io_outAct),
    .io_inwtValid(PEs_4_7_io_inwtValid)
  );
  PE PEs_4_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_8_clock),
    .io_inAct(PEs_4_8_io_inAct),
    .io_inWtPS(PEs_4_8_io_inWtPS),
    .io_outWtPS(PEs_4_8_io_outWtPS),
    .io_outAct(PEs_4_8_io_outAct),
    .io_inwtValid(PEs_4_8_io_inwtValid)
  );
  PE PEs_4_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_9_clock),
    .io_inAct(PEs_4_9_io_inAct),
    .io_inWtPS(PEs_4_9_io_inWtPS),
    .io_outWtPS(PEs_4_9_io_outWtPS),
    .io_outAct(PEs_4_9_io_outAct),
    .io_inwtValid(PEs_4_9_io_inwtValid)
  );
  PE PEs_5_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_0_clock),
    .io_inAct(PEs_5_0_io_inAct),
    .io_inWtPS(PEs_5_0_io_inWtPS),
    .io_outWtPS(PEs_5_0_io_outWtPS),
    .io_outAct(PEs_5_0_io_outAct),
    .io_inwtValid(PEs_5_0_io_inwtValid)
  );
  PE PEs_5_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_1_clock),
    .io_inAct(PEs_5_1_io_inAct),
    .io_inWtPS(PEs_5_1_io_inWtPS),
    .io_outWtPS(PEs_5_1_io_outWtPS),
    .io_outAct(PEs_5_1_io_outAct),
    .io_inwtValid(PEs_5_1_io_inwtValid)
  );
  PE PEs_5_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_2_clock),
    .io_inAct(PEs_5_2_io_inAct),
    .io_inWtPS(PEs_5_2_io_inWtPS),
    .io_outWtPS(PEs_5_2_io_outWtPS),
    .io_outAct(PEs_5_2_io_outAct),
    .io_inwtValid(PEs_5_2_io_inwtValid)
  );
  PE PEs_5_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_3_clock),
    .io_inAct(PEs_5_3_io_inAct),
    .io_inWtPS(PEs_5_3_io_inWtPS),
    .io_outWtPS(PEs_5_3_io_outWtPS),
    .io_outAct(PEs_5_3_io_outAct),
    .io_inwtValid(PEs_5_3_io_inwtValid)
  );
  PE PEs_5_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_4_clock),
    .io_inAct(PEs_5_4_io_inAct),
    .io_inWtPS(PEs_5_4_io_inWtPS),
    .io_outWtPS(PEs_5_4_io_outWtPS),
    .io_outAct(PEs_5_4_io_outAct),
    .io_inwtValid(PEs_5_4_io_inwtValid)
  );
  PE PEs_5_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_5_clock),
    .io_inAct(PEs_5_5_io_inAct),
    .io_inWtPS(PEs_5_5_io_inWtPS),
    .io_outWtPS(PEs_5_5_io_outWtPS),
    .io_outAct(PEs_5_5_io_outAct),
    .io_inwtValid(PEs_5_5_io_inwtValid)
  );
  PE PEs_5_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_6_clock),
    .io_inAct(PEs_5_6_io_inAct),
    .io_inWtPS(PEs_5_6_io_inWtPS),
    .io_outWtPS(PEs_5_6_io_outWtPS),
    .io_outAct(PEs_5_6_io_outAct),
    .io_inwtValid(PEs_5_6_io_inwtValid)
  );
  PE PEs_5_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_7_clock),
    .io_inAct(PEs_5_7_io_inAct),
    .io_inWtPS(PEs_5_7_io_inWtPS),
    .io_outWtPS(PEs_5_7_io_outWtPS),
    .io_outAct(PEs_5_7_io_outAct),
    .io_inwtValid(PEs_5_7_io_inwtValid)
  );
  PE PEs_5_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_8_clock),
    .io_inAct(PEs_5_8_io_inAct),
    .io_inWtPS(PEs_5_8_io_inWtPS),
    .io_outWtPS(PEs_5_8_io_outWtPS),
    .io_outAct(PEs_5_8_io_outAct),
    .io_inwtValid(PEs_5_8_io_inwtValid)
  );
  PE PEs_5_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_9_clock),
    .io_inAct(PEs_5_9_io_inAct),
    .io_inWtPS(PEs_5_9_io_inWtPS),
    .io_outWtPS(PEs_5_9_io_outWtPS),
    .io_outAct(PEs_5_9_io_outAct),
    .io_inwtValid(PEs_5_9_io_inwtValid)
  );
  PE PEs_6_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_0_clock),
    .io_inAct(PEs_6_0_io_inAct),
    .io_inWtPS(PEs_6_0_io_inWtPS),
    .io_outWtPS(PEs_6_0_io_outWtPS),
    .io_outAct(PEs_6_0_io_outAct),
    .io_inwtValid(PEs_6_0_io_inwtValid)
  );
  PE PEs_6_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_1_clock),
    .io_inAct(PEs_6_1_io_inAct),
    .io_inWtPS(PEs_6_1_io_inWtPS),
    .io_outWtPS(PEs_6_1_io_outWtPS),
    .io_outAct(PEs_6_1_io_outAct),
    .io_inwtValid(PEs_6_1_io_inwtValid)
  );
  PE PEs_6_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_2_clock),
    .io_inAct(PEs_6_2_io_inAct),
    .io_inWtPS(PEs_6_2_io_inWtPS),
    .io_outWtPS(PEs_6_2_io_outWtPS),
    .io_outAct(PEs_6_2_io_outAct),
    .io_inwtValid(PEs_6_2_io_inwtValid)
  );
  PE PEs_6_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_3_clock),
    .io_inAct(PEs_6_3_io_inAct),
    .io_inWtPS(PEs_6_3_io_inWtPS),
    .io_outWtPS(PEs_6_3_io_outWtPS),
    .io_outAct(PEs_6_3_io_outAct),
    .io_inwtValid(PEs_6_3_io_inwtValid)
  );
  PE PEs_6_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_4_clock),
    .io_inAct(PEs_6_4_io_inAct),
    .io_inWtPS(PEs_6_4_io_inWtPS),
    .io_outWtPS(PEs_6_4_io_outWtPS),
    .io_outAct(PEs_6_4_io_outAct),
    .io_inwtValid(PEs_6_4_io_inwtValid)
  );
  PE PEs_6_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_5_clock),
    .io_inAct(PEs_6_5_io_inAct),
    .io_inWtPS(PEs_6_5_io_inWtPS),
    .io_outWtPS(PEs_6_5_io_outWtPS),
    .io_outAct(PEs_6_5_io_outAct),
    .io_inwtValid(PEs_6_5_io_inwtValid)
  );
  PE PEs_6_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_6_clock),
    .io_inAct(PEs_6_6_io_inAct),
    .io_inWtPS(PEs_6_6_io_inWtPS),
    .io_outWtPS(PEs_6_6_io_outWtPS),
    .io_outAct(PEs_6_6_io_outAct),
    .io_inwtValid(PEs_6_6_io_inwtValid)
  );
  PE PEs_6_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_7_clock),
    .io_inAct(PEs_6_7_io_inAct),
    .io_inWtPS(PEs_6_7_io_inWtPS),
    .io_outWtPS(PEs_6_7_io_outWtPS),
    .io_outAct(PEs_6_7_io_outAct),
    .io_inwtValid(PEs_6_7_io_inwtValid)
  );
  PE PEs_6_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_8_clock),
    .io_inAct(PEs_6_8_io_inAct),
    .io_inWtPS(PEs_6_8_io_inWtPS),
    .io_outWtPS(PEs_6_8_io_outWtPS),
    .io_outAct(PEs_6_8_io_outAct),
    .io_inwtValid(PEs_6_8_io_inwtValid)
  );
  PE PEs_6_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_9_clock),
    .io_inAct(PEs_6_9_io_inAct),
    .io_inWtPS(PEs_6_9_io_inWtPS),
    .io_outWtPS(PEs_6_9_io_outWtPS),
    .io_outAct(PEs_6_9_io_outAct),
    .io_inwtValid(PEs_6_9_io_inwtValid)
  );
  PE PEs_7_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_0_clock),
    .io_inAct(PEs_7_0_io_inAct),
    .io_inWtPS(PEs_7_0_io_inWtPS),
    .io_outWtPS(PEs_7_0_io_outWtPS),
    .io_outAct(PEs_7_0_io_outAct),
    .io_inwtValid(PEs_7_0_io_inwtValid)
  );
  PE PEs_7_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_1_clock),
    .io_inAct(PEs_7_1_io_inAct),
    .io_inWtPS(PEs_7_1_io_inWtPS),
    .io_outWtPS(PEs_7_1_io_outWtPS),
    .io_outAct(PEs_7_1_io_outAct),
    .io_inwtValid(PEs_7_1_io_inwtValid)
  );
  PE PEs_7_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_2_clock),
    .io_inAct(PEs_7_2_io_inAct),
    .io_inWtPS(PEs_7_2_io_inWtPS),
    .io_outWtPS(PEs_7_2_io_outWtPS),
    .io_outAct(PEs_7_2_io_outAct),
    .io_inwtValid(PEs_7_2_io_inwtValid)
  );
  PE PEs_7_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_3_clock),
    .io_inAct(PEs_7_3_io_inAct),
    .io_inWtPS(PEs_7_3_io_inWtPS),
    .io_outWtPS(PEs_7_3_io_outWtPS),
    .io_outAct(PEs_7_3_io_outAct),
    .io_inwtValid(PEs_7_3_io_inwtValid)
  );
  PE PEs_7_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_4_clock),
    .io_inAct(PEs_7_4_io_inAct),
    .io_inWtPS(PEs_7_4_io_inWtPS),
    .io_outWtPS(PEs_7_4_io_outWtPS),
    .io_outAct(PEs_7_4_io_outAct),
    .io_inwtValid(PEs_7_4_io_inwtValid)
  );
  PE PEs_7_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_5_clock),
    .io_inAct(PEs_7_5_io_inAct),
    .io_inWtPS(PEs_7_5_io_inWtPS),
    .io_outWtPS(PEs_7_5_io_outWtPS),
    .io_outAct(PEs_7_5_io_outAct),
    .io_inwtValid(PEs_7_5_io_inwtValid)
  );
  PE PEs_7_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_6_clock),
    .io_inAct(PEs_7_6_io_inAct),
    .io_inWtPS(PEs_7_6_io_inWtPS),
    .io_outWtPS(PEs_7_6_io_outWtPS),
    .io_outAct(PEs_7_6_io_outAct),
    .io_inwtValid(PEs_7_6_io_inwtValid)
  );
  PE PEs_7_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_7_clock),
    .io_inAct(PEs_7_7_io_inAct),
    .io_inWtPS(PEs_7_7_io_inWtPS),
    .io_outWtPS(PEs_7_7_io_outWtPS),
    .io_outAct(PEs_7_7_io_outAct),
    .io_inwtValid(PEs_7_7_io_inwtValid)
  );
  PE PEs_7_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_8_clock),
    .io_inAct(PEs_7_8_io_inAct),
    .io_inWtPS(PEs_7_8_io_inWtPS),
    .io_outWtPS(PEs_7_8_io_outWtPS),
    .io_outAct(PEs_7_8_io_outAct),
    .io_inwtValid(PEs_7_8_io_inwtValid)
  );
  PE PEs_7_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_9_clock),
    .io_inAct(PEs_7_9_io_inAct),
    .io_inWtPS(PEs_7_9_io_inWtPS),
    .io_outWtPS(PEs_7_9_io_outWtPS),
    .io_outAct(PEs_7_9_io_outAct),
    .io_inwtValid(PEs_7_9_io_inwtValid)
  );
  PE PEs_8_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_0_clock),
    .io_inAct(PEs_8_0_io_inAct),
    .io_inWtPS(PEs_8_0_io_inWtPS),
    .io_outWtPS(PEs_8_0_io_outWtPS),
    .io_outAct(PEs_8_0_io_outAct),
    .io_inwtValid(PEs_8_0_io_inwtValid)
  );
  PE PEs_8_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_1_clock),
    .io_inAct(PEs_8_1_io_inAct),
    .io_inWtPS(PEs_8_1_io_inWtPS),
    .io_outWtPS(PEs_8_1_io_outWtPS),
    .io_outAct(PEs_8_1_io_outAct),
    .io_inwtValid(PEs_8_1_io_inwtValid)
  );
  PE PEs_8_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_2_clock),
    .io_inAct(PEs_8_2_io_inAct),
    .io_inWtPS(PEs_8_2_io_inWtPS),
    .io_outWtPS(PEs_8_2_io_outWtPS),
    .io_outAct(PEs_8_2_io_outAct),
    .io_inwtValid(PEs_8_2_io_inwtValid)
  );
  PE PEs_8_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_3_clock),
    .io_inAct(PEs_8_3_io_inAct),
    .io_inWtPS(PEs_8_3_io_inWtPS),
    .io_outWtPS(PEs_8_3_io_outWtPS),
    .io_outAct(PEs_8_3_io_outAct),
    .io_inwtValid(PEs_8_3_io_inwtValid)
  );
  PE PEs_8_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_4_clock),
    .io_inAct(PEs_8_4_io_inAct),
    .io_inWtPS(PEs_8_4_io_inWtPS),
    .io_outWtPS(PEs_8_4_io_outWtPS),
    .io_outAct(PEs_8_4_io_outAct),
    .io_inwtValid(PEs_8_4_io_inwtValid)
  );
  PE PEs_8_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_5_clock),
    .io_inAct(PEs_8_5_io_inAct),
    .io_inWtPS(PEs_8_5_io_inWtPS),
    .io_outWtPS(PEs_8_5_io_outWtPS),
    .io_outAct(PEs_8_5_io_outAct),
    .io_inwtValid(PEs_8_5_io_inwtValid)
  );
  PE PEs_8_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_6_clock),
    .io_inAct(PEs_8_6_io_inAct),
    .io_inWtPS(PEs_8_6_io_inWtPS),
    .io_outWtPS(PEs_8_6_io_outWtPS),
    .io_outAct(PEs_8_6_io_outAct),
    .io_inwtValid(PEs_8_6_io_inwtValid)
  );
  PE PEs_8_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_7_clock),
    .io_inAct(PEs_8_7_io_inAct),
    .io_inWtPS(PEs_8_7_io_inWtPS),
    .io_outWtPS(PEs_8_7_io_outWtPS),
    .io_outAct(PEs_8_7_io_outAct),
    .io_inwtValid(PEs_8_7_io_inwtValid)
  );
  PE PEs_8_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_8_clock),
    .io_inAct(PEs_8_8_io_inAct),
    .io_inWtPS(PEs_8_8_io_inWtPS),
    .io_outWtPS(PEs_8_8_io_outWtPS),
    .io_outAct(PEs_8_8_io_outAct),
    .io_inwtValid(PEs_8_8_io_inwtValid)
  );
  PE PEs_8_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_9_clock),
    .io_inAct(PEs_8_9_io_inAct),
    .io_inWtPS(PEs_8_9_io_inWtPS),
    .io_outWtPS(PEs_8_9_io_outWtPS),
    .io_outAct(PEs_8_9_io_outAct),
    .io_inwtValid(PEs_8_9_io_inwtValid)
  );
  PE PEs_9_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_0_clock),
    .io_inAct(PEs_9_0_io_inAct),
    .io_inWtPS(PEs_9_0_io_inWtPS),
    .io_outWtPS(PEs_9_0_io_outWtPS),
    .io_outAct(PEs_9_0_io_outAct),
    .io_inwtValid(PEs_9_0_io_inwtValid)
  );
  PE PEs_9_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_1_clock),
    .io_inAct(PEs_9_1_io_inAct),
    .io_inWtPS(PEs_9_1_io_inWtPS),
    .io_outWtPS(PEs_9_1_io_outWtPS),
    .io_outAct(PEs_9_1_io_outAct),
    .io_inwtValid(PEs_9_1_io_inwtValid)
  );
  PE PEs_9_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_2_clock),
    .io_inAct(PEs_9_2_io_inAct),
    .io_inWtPS(PEs_9_2_io_inWtPS),
    .io_outWtPS(PEs_9_2_io_outWtPS),
    .io_outAct(PEs_9_2_io_outAct),
    .io_inwtValid(PEs_9_2_io_inwtValid)
  );
  PE PEs_9_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_3_clock),
    .io_inAct(PEs_9_3_io_inAct),
    .io_inWtPS(PEs_9_3_io_inWtPS),
    .io_outWtPS(PEs_9_3_io_outWtPS),
    .io_outAct(PEs_9_3_io_outAct),
    .io_inwtValid(PEs_9_3_io_inwtValid)
  );
  PE PEs_9_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_4_clock),
    .io_inAct(PEs_9_4_io_inAct),
    .io_inWtPS(PEs_9_4_io_inWtPS),
    .io_outWtPS(PEs_9_4_io_outWtPS),
    .io_outAct(PEs_9_4_io_outAct),
    .io_inwtValid(PEs_9_4_io_inwtValid)
  );
  PE PEs_9_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_5_clock),
    .io_inAct(PEs_9_5_io_inAct),
    .io_inWtPS(PEs_9_5_io_inWtPS),
    .io_outWtPS(PEs_9_5_io_outWtPS),
    .io_outAct(PEs_9_5_io_outAct),
    .io_inwtValid(PEs_9_5_io_inwtValid)
  );
  PE PEs_9_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_6_clock),
    .io_inAct(PEs_9_6_io_inAct),
    .io_inWtPS(PEs_9_6_io_inWtPS),
    .io_outWtPS(PEs_9_6_io_outWtPS),
    .io_outAct(PEs_9_6_io_outAct),
    .io_inwtValid(PEs_9_6_io_inwtValid)
  );
  PE PEs_9_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_7_clock),
    .io_inAct(PEs_9_7_io_inAct),
    .io_inWtPS(PEs_9_7_io_inWtPS),
    .io_outWtPS(PEs_9_7_io_outWtPS),
    .io_outAct(PEs_9_7_io_outAct),
    .io_inwtValid(PEs_9_7_io_inwtValid)
  );
  PE PEs_9_8 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_8_clock),
    .io_inAct(PEs_9_8_io_inAct),
    .io_inWtPS(PEs_9_8_io_inWtPS),
    .io_outWtPS(PEs_9_8_io_outWtPS),
    .io_outAct(PEs_9_8_io_outAct),
    .io_inwtValid(PEs_9_8_io_inwtValid)
  );
  PE PEs_9_9 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_9_clock),
    .io_inAct(PEs_9_9_io_inAct),
    .io_inWtPS(PEs_9_9_io_inWtPS),
    .io_outWtPS(PEs_9_9_io_outWtPS),
    .io_outAct(PEs_9_9_io_outAct),
    .io_inwtValid(PEs_9_9_io_inwtValid)
  );
  assign io_outSum_0 = PEs_9_0_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_1 = PEs_9_1_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_2 = PEs_9_2_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_3 = PEs_9_3_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_4 = PEs_9_4_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_5 = PEs_9_5_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_6 = PEs_9_6_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_7 = PEs_9_7_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_8 = PEs_9_8_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_9 = PEs_9_9_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign PEs_0_0_clock = clock;
  assign PEs_0_0_io_inAct = io_inAct_0; // @[SystolicArray.scala 38:44]
  assign PEs_0_0_io_inWtPS = {{24{io_inWeight_0[15]}},io_inWeight_0}; // @[SystolicArray.scala 31:45]
  assign PEs_0_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_1_clock = clock;
  assign PEs_0_1_io_inAct = PEs_0_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_1_io_inWtPS = {{24{io_inWeight_1[15]}},io_inWeight_1}; // @[SystolicArray.scala 31:45]
  assign PEs_0_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_2_clock = clock;
  assign PEs_0_2_io_inAct = PEs_0_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_2_io_inWtPS = {{24{io_inWeight_2[15]}},io_inWeight_2}; // @[SystolicArray.scala 31:45]
  assign PEs_0_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_3_clock = clock;
  assign PEs_0_3_io_inAct = PEs_0_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_3_io_inWtPS = {{24{io_inWeight_3[15]}},io_inWeight_3}; // @[SystolicArray.scala 31:45]
  assign PEs_0_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_4_clock = clock;
  assign PEs_0_4_io_inAct = PEs_0_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_4_io_inWtPS = {{24{io_inWeight_4[15]}},io_inWeight_4}; // @[SystolicArray.scala 31:45]
  assign PEs_0_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_5_clock = clock;
  assign PEs_0_5_io_inAct = PEs_0_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_5_io_inWtPS = {{24{io_inWeight_5[15]}},io_inWeight_5}; // @[SystolicArray.scala 31:45]
  assign PEs_0_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_6_clock = clock;
  assign PEs_0_6_io_inAct = PEs_0_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_6_io_inWtPS = {{24{io_inWeight_6[15]}},io_inWeight_6}; // @[SystolicArray.scala 31:45]
  assign PEs_0_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_7_clock = clock;
  assign PEs_0_7_io_inAct = PEs_0_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_7_io_inWtPS = {{24{io_inWeight_7[15]}},io_inWeight_7}; // @[SystolicArray.scala 31:45]
  assign PEs_0_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_8_clock = clock;
  assign PEs_0_8_io_inAct = PEs_0_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_8_io_inWtPS = {{24{io_inWeight_8[15]}},io_inWeight_8}; // @[SystolicArray.scala 31:45]
  assign PEs_0_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_9_clock = clock;
  assign PEs_0_9_io_inAct = PEs_0_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_9_io_inWtPS = {{24{io_inWeight_9[15]}},io_inWeight_9}; // @[SystolicArray.scala 31:45]
  assign PEs_0_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_0_clock = clock;
  assign PEs_1_0_io_inAct = io_inAct_1; // @[SystolicArray.scala 38:44]
  assign PEs_1_0_io_inWtPS = PEs_0_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_1_clock = clock;
  assign PEs_1_1_io_inAct = PEs_1_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_1_io_inWtPS = PEs_0_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_2_clock = clock;
  assign PEs_1_2_io_inAct = PEs_1_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_2_io_inWtPS = PEs_0_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_3_clock = clock;
  assign PEs_1_3_io_inAct = PEs_1_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_3_io_inWtPS = PEs_0_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_4_clock = clock;
  assign PEs_1_4_io_inAct = PEs_1_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_4_io_inWtPS = PEs_0_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_5_clock = clock;
  assign PEs_1_5_io_inAct = PEs_1_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_5_io_inWtPS = PEs_0_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_6_clock = clock;
  assign PEs_1_6_io_inAct = PEs_1_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_6_io_inWtPS = PEs_0_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_7_clock = clock;
  assign PEs_1_7_io_inAct = PEs_1_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_7_io_inWtPS = PEs_0_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_8_clock = clock;
  assign PEs_1_8_io_inAct = PEs_1_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_8_io_inWtPS = PEs_0_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_9_clock = clock;
  assign PEs_1_9_io_inAct = PEs_1_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_9_io_inWtPS = PEs_0_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_0_clock = clock;
  assign PEs_2_0_io_inAct = io_inAct_2; // @[SystolicArray.scala 38:44]
  assign PEs_2_0_io_inWtPS = PEs_1_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_1_clock = clock;
  assign PEs_2_1_io_inAct = PEs_2_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_1_io_inWtPS = PEs_1_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_2_clock = clock;
  assign PEs_2_2_io_inAct = PEs_2_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_2_io_inWtPS = PEs_1_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_3_clock = clock;
  assign PEs_2_3_io_inAct = PEs_2_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_3_io_inWtPS = PEs_1_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_4_clock = clock;
  assign PEs_2_4_io_inAct = PEs_2_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_4_io_inWtPS = PEs_1_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_5_clock = clock;
  assign PEs_2_5_io_inAct = PEs_2_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_5_io_inWtPS = PEs_1_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_6_clock = clock;
  assign PEs_2_6_io_inAct = PEs_2_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_6_io_inWtPS = PEs_1_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_7_clock = clock;
  assign PEs_2_7_io_inAct = PEs_2_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_7_io_inWtPS = PEs_1_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_8_clock = clock;
  assign PEs_2_8_io_inAct = PEs_2_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_8_io_inWtPS = PEs_1_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_9_clock = clock;
  assign PEs_2_9_io_inAct = PEs_2_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_9_io_inWtPS = PEs_1_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_0_clock = clock;
  assign PEs_3_0_io_inAct = io_inAct_3; // @[SystolicArray.scala 38:44]
  assign PEs_3_0_io_inWtPS = PEs_2_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_1_clock = clock;
  assign PEs_3_1_io_inAct = PEs_3_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_1_io_inWtPS = PEs_2_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_2_clock = clock;
  assign PEs_3_2_io_inAct = PEs_3_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_2_io_inWtPS = PEs_2_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_3_clock = clock;
  assign PEs_3_3_io_inAct = PEs_3_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_3_io_inWtPS = PEs_2_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_4_clock = clock;
  assign PEs_3_4_io_inAct = PEs_3_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_4_io_inWtPS = PEs_2_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_5_clock = clock;
  assign PEs_3_5_io_inAct = PEs_3_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_5_io_inWtPS = PEs_2_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_6_clock = clock;
  assign PEs_3_6_io_inAct = PEs_3_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_6_io_inWtPS = PEs_2_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_7_clock = clock;
  assign PEs_3_7_io_inAct = PEs_3_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_7_io_inWtPS = PEs_2_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_8_clock = clock;
  assign PEs_3_8_io_inAct = PEs_3_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_8_io_inWtPS = PEs_2_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_9_clock = clock;
  assign PEs_3_9_io_inAct = PEs_3_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_9_io_inWtPS = PEs_2_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_0_clock = clock;
  assign PEs_4_0_io_inAct = io_inAct_4; // @[SystolicArray.scala 38:44]
  assign PEs_4_0_io_inWtPS = PEs_3_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_1_clock = clock;
  assign PEs_4_1_io_inAct = PEs_4_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_1_io_inWtPS = PEs_3_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_2_clock = clock;
  assign PEs_4_2_io_inAct = PEs_4_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_2_io_inWtPS = PEs_3_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_3_clock = clock;
  assign PEs_4_3_io_inAct = PEs_4_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_3_io_inWtPS = PEs_3_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_4_clock = clock;
  assign PEs_4_4_io_inAct = PEs_4_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_4_io_inWtPS = PEs_3_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_5_clock = clock;
  assign PEs_4_5_io_inAct = PEs_4_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_5_io_inWtPS = PEs_3_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_6_clock = clock;
  assign PEs_4_6_io_inAct = PEs_4_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_6_io_inWtPS = PEs_3_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_7_clock = clock;
  assign PEs_4_7_io_inAct = PEs_4_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_7_io_inWtPS = PEs_3_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_8_clock = clock;
  assign PEs_4_8_io_inAct = PEs_4_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_8_io_inWtPS = PEs_3_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_9_clock = clock;
  assign PEs_4_9_io_inAct = PEs_4_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_9_io_inWtPS = PEs_3_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_0_clock = clock;
  assign PEs_5_0_io_inAct = io_inAct_5; // @[SystolicArray.scala 38:44]
  assign PEs_5_0_io_inWtPS = PEs_4_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_1_clock = clock;
  assign PEs_5_1_io_inAct = PEs_5_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_1_io_inWtPS = PEs_4_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_2_clock = clock;
  assign PEs_5_2_io_inAct = PEs_5_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_2_io_inWtPS = PEs_4_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_3_clock = clock;
  assign PEs_5_3_io_inAct = PEs_5_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_3_io_inWtPS = PEs_4_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_4_clock = clock;
  assign PEs_5_4_io_inAct = PEs_5_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_4_io_inWtPS = PEs_4_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_5_clock = clock;
  assign PEs_5_5_io_inAct = PEs_5_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_5_io_inWtPS = PEs_4_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_6_clock = clock;
  assign PEs_5_6_io_inAct = PEs_5_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_6_io_inWtPS = PEs_4_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_7_clock = clock;
  assign PEs_5_7_io_inAct = PEs_5_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_7_io_inWtPS = PEs_4_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_8_clock = clock;
  assign PEs_5_8_io_inAct = PEs_5_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_8_io_inWtPS = PEs_4_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_9_clock = clock;
  assign PEs_5_9_io_inAct = PEs_5_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_9_io_inWtPS = PEs_4_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_0_clock = clock;
  assign PEs_6_0_io_inAct = io_inAct_6; // @[SystolicArray.scala 38:44]
  assign PEs_6_0_io_inWtPS = PEs_5_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_1_clock = clock;
  assign PEs_6_1_io_inAct = PEs_6_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_1_io_inWtPS = PEs_5_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_2_clock = clock;
  assign PEs_6_2_io_inAct = PEs_6_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_2_io_inWtPS = PEs_5_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_3_clock = clock;
  assign PEs_6_3_io_inAct = PEs_6_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_3_io_inWtPS = PEs_5_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_4_clock = clock;
  assign PEs_6_4_io_inAct = PEs_6_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_4_io_inWtPS = PEs_5_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_5_clock = clock;
  assign PEs_6_5_io_inAct = PEs_6_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_5_io_inWtPS = PEs_5_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_6_clock = clock;
  assign PEs_6_6_io_inAct = PEs_6_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_6_io_inWtPS = PEs_5_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_7_clock = clock;
  assign PEs_6_7_io_inAct = PEs_6_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_7_io_inWtPS = PEs_5_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_8_clock = clock;
  assign PEs_6_8_io_inAct = PEs_6_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_8_io_inWtPS = PEs_5_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_9_clock = clock;
  assign PEs_6_9_io_inAct = PEs_6_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_9_io_inWtPS = PEs_5_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_0_clock = clock;
  assign PEs_7_0_io_inAct = io_inAct_7; // @[SystolicArray.scala 38:44]
  assign PEs_7_0_io_inWtPS = PEs_6_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_1_clock = clock;
  assign PEs_7_1_io_inAct = PEs_7_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_1_io_inWtPS = PEs_6_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_2_clock = clock;
  assign PEs_7_2_io_inAct = PEs_7_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_2_io_inWtPS = PEs_6_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_3_clock = clock;
  assign PEs_7_3_io_inAct = PEs_7_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_3_io_inWtPS = PEs_6_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_4_clock = clock;
  assign PEs_7_4_io_inAct = PEs_7_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_4_io_inWtPS = PEs_6_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_5_clock = clock;
  assign PEs_7_5_io_inAct = PEs_7_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_5_io_inWtPS = PEs_6_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_6_clock = clock;
  assign PEs_7_6_io_inAct = PEs_7_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_6_io_inWtPS = PEs_6_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_7_clock = clock;
  assign PEs_7_7_io_inAct = PEs_7_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_7_io_inWtPS = PEs_6_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_8_clock = clock;
  assign PEs_7_8_io_inAct = PEs_7_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_8_io_inWtPS = PEs_6_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_9_clock = clock;
  assign PEs_7_9_io_inAct = PEs_7_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_9_io_inWtPS = PEs_6_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_0_clock = clock;
  assign PEs_8_0_io_inAct = io_inAct_8; // @[SystolicArray.scala 38:44]
  assign PEs_8_0_io_inWtPS = PEs_7_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_1_clock = clock;
  assign PEs_8_1_io_inAct = PEs_8_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_1_io_inWtPS = PEs_7_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_2_clock = clock;
  assign PEs_8_2_io_inAct = PEs_8_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_2_io_inWtPS = PEs_7_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_3_clock = clock;
  assign PEs_8_3_io_inAct = PEs_8_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_3_io_inWtPS = PEs_7_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_4_clock = clock;
  assign PEs_8_4_io_inAct = PEs_8_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_4_io_inWtPS = PEs_7_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_5_clock = clock;
  assign PEs_8_5_io_inAct = PEs_8_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_5_io_inWtPS = PEs_7_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_6_clock = clock;
  assign PEs_8_6_io_inAct = PEs_8_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_6_io_inWtPS = PEs_7_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_7_clock = clock;
  assign PEs_8_7_io_inAct = PEs_8_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_7_io_inWtPS = PEs_7_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_8_clock = clock;
  assign PEs_8_8_io_inAct = PEs_8_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_8_io_inWtPS = PEs_7_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_9_clock = clock;
  assign PEs_8_9_io_inAct = PEs_8_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_9_io_inWtPS = PEs_7_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_0_clock = clock;
  assign PEs_9_0_io_inAct = io_inAct_9; // @[SystolicArray.scala 38:44]
  assign PEs_9_0_io_inWtPS = PEs_8_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_1_clock = clock;
  assign PEs_9_1_io_inAct = PEs_9_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_1_io_inWtPS = PEs_8_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_2_clock = clock;
  assign PEs_9_2_io_inAct = PEs_9_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_2_io_inWtPS = PEs_8_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_3_clock = clock;
  assign PEs_9_3_io_inAct = PEs_9_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_3_io_inWtPS = PEs_8_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_4_clock = clock;
  assign PEs_9_4_io_inAct = PEs_9_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_4_io_inWtPS = PEs_8_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_5_clock = clock;
  assign PEs_9_5_io_inAct = PEs_9_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_5_io_inWtPS = PEs_8_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_6_clock = clock;
  assign PEs_9_6_io_inAct = PEs_9_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_6_io_inWtPS = PEs_8_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_7_clock = clock;
  assign PEs_9_7_io_inAct = PEs_9_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_7_io_inWtPS = PEs_8_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_8_clock = clock;
  assign PEs_9_8_io_inAct = PEs_9_7_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_8_io_inWtPS = PEs_8_8_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_8_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_9_clock = clock;
  assign PEs_9_9_io_inAct = PEs_9_8_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_9_io_inWtPS = PEs_8_9_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_9_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  always @(posedge clock) begin
    validReg <= io_inwtValid; // @[SystolicArray.scala 22:25]
  end
endmodule
module SystolicArray_2(
  input         clock,
  input  [15:0] io_inAct_0,
  input  [15:0] io_inAct_1,
  input  [15:0] io_inAct_2,
  input  [15:0] io_inAct_3,
  input  [15:0] io_inAct_4,
  input  [15:0] io_inAct_5,
  input  [15:0] io_inAct_6,
  input  [15:0] io_inAct_7,
  input  [15:0] io_inAct_8,
  input  [15:0] io_inAct_9,
  input  [15:0] io_inWeight_0,
  input  [15:0] io_inWeight_1,
  input  [15:0] io_inWeight_2,
  input  [15:0] io_inWeight_3,
  input  [15:0] io_inWeight_4,
  input  [15:0] io_inWeight_5,
  input  [15:0] io_inWeight_6,
  input  [15:0] io_inWeight_7,
  output [39:0] io_outSum_0,
  output [39:0] io_outSum_1,
  output [39:0] io_outSum_2,
  output [39:0] io_outSum_3,
  output [39:0] io_outSum_4,
  output [39:0] io_outSum_5,
  output [39:0] io_outSum_6,
  output [39:0] io_outSum_7,
  input         io_inwtValid
);
  wire  PEs_0_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_0_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_0_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_0_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_1_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_1_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_1_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_2_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_2_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_2_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_3_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_3_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_3_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_4_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_4_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_4_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_5_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_5_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_5_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_6_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_6_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_6_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_7_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_7_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_7_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_8_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_8_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_8_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_0_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_0_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_0_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_1_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_1_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_1_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_2_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_2_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_2_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_3_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_3_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_3_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_4_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_4_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_4_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_5_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_5_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_5_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_6_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_6_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_6_io_inwtValid; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_clock; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_inAct; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_inWtPS; // @[SystolicArray.scala 18:65]
  wire [39:0] PEs_9_7_io_outWtPS; // @[SystolicArray.scala 18:65]
  wire [15:0] PEs_9_7_io_outAct; // @[SystolicArray.scala 18:65]
  wire  PEs_9_7_io_inwtValid; // @[SystolicArray.scala 18:65]
  reg  validReg; // @[SystolicArray.scala 22:25]
  PE PEs_0_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_0_clock),
    .io_inAct(PEs_0_0_io_inAct),
    .io_inWtPS(PEs_0_0_io_inWtPS),
    .io_outWtPS(PEs_0_0_io_outWtPS),
    .io_outAct(PEs_0_0_io_outAct),
    .io_inwtValid(PEs_0_0_io_inwtValid)
  );
  PE PEs_0_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_1_clock),
    .io_inAct(PEs_0_1_io_inAct),
    .io_inWtPS(PEs_0_1_io_inWtPS),
    .io_outWtPS(PEs_0_1_io_outWtPS),
    .io_outAct(PEs_0_1_io_outAct),
    .io_inwtValid(PEs_0_1_io_inwtValid)
  );
  PE PEs_0_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_2_clock),
    .io_inAct(PEs_0_2_io_inAct),
    .io_inWtPS(PEs_0_2_io_inWtPS),
    .io_outWtPS(PEs_0_2_io_outWtPS),
    .io_outAct(PEs_0_2_io_outAct),
    .io_inwtValid(PEs_0_2_io_inwtValid)
  );
  PE PEs_0_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_3_clock),
    .io_inAct(PEs_0_3_io_inAct),
    .io_inWtPS(PEs_0_3_io_inWtPS),
    .io_outWtPS(PEs_0_3_io_outWtPS),
    .io_outAct(PEs_0_3_io_outAct),
    .io_inwtValid(PEs_0_3_io_inwtValid)
  );
  PE PEs_0_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_4_clock),
    .io_inAct(PEs_0_4_io_inAct),
    .io_inWtPS(PEs_0_4_io_inWtPS),
    .io_outWtPS(PEs_0_4_io_outWtPS),
    .io_outAct(PEs_0_4_io_outAct),
    .io_inwtValid(PEs_0_4_io_inwtValid)
  );
  PE PEs_0_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_5_clock),
    .io_inAct(PEs_0_5_io_inAct),
    .io_inWtPS(PEs_0_5_io_inWtPS),
    .io_outWtPS(PEs_0_5_io_outWtPS),
    .io_outAct(PEs_0_5_io_outAct),
    .io_inwtValid(PEs_0_5_io_inwtValid)
  );
  PE PEs_0_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_6_clock),
    .io_inAct(PEs_0_6_io_inAct),
    .io_inWtPS(PEs_0_6_io_inWtPS),
    .io_outWtPS(PEs_0_6_io_outWtPS),
    .io_outAct(PEs_0_6_io_outAct),
    .io_inwtValid(PEs_0_6_io_inwtValid)
  );
  PE PEs_0_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_0_7_clock),
    .io_inAct(PEs_0_7_io_inAct),
    .io_inWtPS(PEs_0_7_io_inWtPS),
    .io_outWtPS(PEs_0_7_io_outWtPS),
    .io_outAct(PEs_0_7_io_outAct),
    .io_inwtValid(PEs_0_7_io_inwtValid)
  );
  PE PEs_1_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_0_clock),
    .io_inAct(PEs_1_0_io_inAct),
    .io_inWtPS(PEs_1_0_io_inWtPS),
    .io_outWtPS(PEs_1_0_io_outWtPS),
    .io_outAct(PEs_1_0_io_outAct),
    .io_inwtValid(PEs_1_0_io_inwtValid)
  );
  PE PEs_1_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_1_clock),
    .io_inAct(PEs_1_1_io_inAct),
    .io_inWtPS(PEs_1_1_io_inWtPS),
    .io_outWtPS(PEs_1_1_io_outWtPS),
    .io_outAct(PEs_1_1_io_outAct),
    .io_inwtValid(PEs_1_1_io_inwtValid)
  );
  PE PEs_1_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_2_clock),
    .io_inAct(PEs_1_2_io_inAct),
    .io_inWtPS(PEs_1_2_io_inWtPS),
    .io_outWtPS(PEs_1_2_io_outWtPS),
    .io_outAct(PEs_1_2_io_outAct),
    .io_inwtValid(PEs_1_2_io_inwtValid)
  );
  PE PEs_1_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_3_clock),
    .io_inAct(PEs_1_3_io_inAct),
    .io_inWtPS(PEs_1_3_io_inWtPS),
    .io_outWtPS(PEs_1_3_io_outWtPS),
    .io_outAct(PEs_1_3_io_outAct),
    .io_inwtValid(PEs_1_3_io_inwtValid)
  );
  PE PEs_1_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_4_clock),
    .io_inAct(PEs_1_4_io_inAct),
    .io_inWtPS(PEs_1_4_io_inWtPS),
    .io_outWtPS(PEs_1_4_io_outWtPS),
    .io_outAct(PEs_1_4_io_outAct),
    .io_inwtValid(PEs_1_4_io_inwtValid)
  );
  PE PEs_1_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_5_clock),
    .io_inAct(PEs_1_5_io_inAct),
    .io_inWtPS(PEs_1_5_io_inWtPS),
    .io_outWtPS(PEs_1_5_io_outWtPS),
    .io_outAct(PEs_1_5_io_outAct),
    .io_inwtValid(PEs_1_5_io_inwtValid)
  );
  PE PEs_1_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_6_clock),
    .io_inAct(PEs_1_6_io_inAct),
    .io_inWtPS(PEs_1_6_io_inWtPS),
    .io_outWtPS(PEs_1_6_io_outWtPS),
    .io_outAct(PEs_1_6_io_outAct),
    .io_inwtValid(PEs_1_6_io_inwtValid)
  );
  PE PEs_1_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_1_7_clock),
    .io_inAct(PEs_1_7_io_inAct),
    .io_inWtPS(PEs_1_7_io_inWtPS),
    .io_outWtPS(PEs_1_7_io_outWtPS),
    .io_outAct(PEs_1_7_io_outAct),
    .io_inwtValid(PEs_1_7_io_inwtValid)
  );
  PE PEs_2_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_0_clock),
    .io_inAct(PEs_2_0_io_inAct),
    .io_inWtPS(PEs_2_0_io_inWtPS),
    .io_outWtPS(PEs_2_0_io_outWtPS),
    .io_outAct(PEs_2_0_io_outAct),
    .io_inwtValid(PEs_2_0_io_inwtValid)
  );
  PE PEs_2_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_1_clock),
    .io_inAct(PEs_2_1_io_inAct),
    .io_inWtPS(PEs_2_1_io_inWtPS),
    .io_outWtPS(PEs_2_1_io_outWtPS),
    .io_outAct(PEs_2_1_io_outAct),
    .io_inwtValid(PEs_2_1_io_inwtValid)
  );
  PE PEs_2_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_2_clock),
    .io_inAct(PEs_2_2_io_inAct),
    .io_inWtPS(PEs_2_2_io_inWtPS),
    .io_outWtPS(PEs_2_2_io_outWtPS),
    .io_outAct(PEs_2_2_io_outAct),
    .io_inwtValid(PEs_2_2_io_inwtValid)
  );
  PE PEs_2_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_3_clock),
    .io_inAct(PEs_2_3_io_inAct),
    .io_inWtPS(PEs_2_3_io_inWtPS),
    .io_outWtPS(PEs_2_3_io_outWtPS),
    .io_outAct(PEs_2_3_io_outAct),
    .io_inwtValid(PEs_2_3_io_inwtValid)
  );
  PE PEs_2_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_4_clock),
    .io_inAct(PEs_2_4_io_inAct),
    .io_inWtPS(PEs_2_4_io_inWtPS),
    .io_outWtPS(PEs_2_4_io_outWtPS),
    .io_outAct(PEs_2_4_io_outAct),
    .io_inwtValid(PEs_2_4_io_inwtValid)
  );
  PE PEs_2_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_5_clock),
    .io_inAct(PEs_2_5_io_inAct),
    .io_inWtPS(PEs_2_5_io_inWtPS),
    .io_outWtPS(PEs_2_5_io_outWtPS),
    .io_outAct(PEs_2_5_io_outAct),
    .io_inwtValid(PEs_2_5_io_inwtValid)
  );
  PE PEs_2_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_6_clock),
    .io_inAct(PEs_2_6_io_inAct),
    .io_inWtPS(PEs_2_6_io_inWtPS),
    .io_outWtPS(PEs_2_6_io_outWtPS),
    .io_outAct(PEs_2_6_io_outAct),
    .io_inwtValid(PEs_2_6_io_inwtValid)
  );
  PE PEs_2_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_2_7_clock),
    .io_inAct(PEs_2_7_io_inAct),
    .io_inWtPS(PEs_2_7_io_inWtPS),
    .io_outWtPS(PEs_2_7_io_outWtPS),
    .io_outAct(PEs_2_7_io_outAct),
    .io_inwtValid(PEs_2_7_io_inwtValid)
  );
  PE PEs_3_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_0_clock),
    .io_inAct(PEs_3_0_io_inAct),
    .io_inWtPS(PEs_3_0_io_inWtPS),
    .io_outWtPS(PEs_3_0_io_outWtPS),
    .io_outAct(PEs_3_0_io_outAct),
    .io_inwtValid(PEs_3_0_io_inwtValid)
  );
  PE PEs_3_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_1_clock),
    .io_inAct(PEs_3_1_io_inAct),
    .io_inWtPS(PEs_3_1_io_inWtPS),
    .io_outWtPS(PEs_3_1_io_outWtPS),
    .io_outAct(PEs_3_1_io_outAct),
    .io_inwtValid(PEs_3_1_io_inwtValid)
  );
  PE PEs_3_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_2_clock),
    .io_inAct(PEs_3_2_io_inAct),
    .io_inWtPS(PEs_3_2_io_inWtPS),
    .io_outWtPS(PEs_3_2_io_outWtPS),
    .io_outAct(PEs_3_2_io_outAct),
    .io_inwtValid(PEs_3_2_io_inwtValid)
  );
  PE PEs_3_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_3_clock),
    .io_inAct(PEs_3_3_io_inAct),
    .io_inWtPS(PEs_3_3_io_inWtPS),
    .io_outWtPS(PEs_3_3_io_outWtPS),
    .io_outAct(PEs_3_3_io_outAct),
    .io_inwtValid(PEs_3_3_io_inwtValid)
  );
  PE PEs_3_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_4_clock),
    .io_inAct(PEs_3_4_io_inAct),
    .io_inWtPS(PEs_3_4_io_inWtPS),
    .io_outWtPS(PEs_3_4_io_outWtPS),
    .io_outAct(PEs_3_4_io_outAct),
    .io_inwtValid(PEs_3_4_io_inwtValid)
  );
  PE PEs_3_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_5_clock),
    .io_inAct(PEs_3_5_io_inAct),
    .io_inWtPS(PEs_3_5_io_inWtPS),
    .io_outWtPS(PEs_3_5_io_outWtPS),
    .io_outAct(PEs_3_5_io_outAct),
    .io_inwtValid(PEs_3_5_io_inwtValid)
  );
  PE PEs_3_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_6_clock),
    .io_inAct(PEs_3_6_io_inAct),
    .io_inWtPS(PEs_3_6_io_inWtPS),
    .io_outWtPS(PEs_3_6_io_outWtPS),
    .io_outAct(PEs_3_6_io_outAct),
    .io_inwtValid(PEs_3_6_io_inwtValid)
  );
  PE PEs_3_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_3_7_clock),
    .io_inAct(PEs_3_7_io_inAct),
    .io_inWtPS(PEs_3_7_io_inWtPS),
    .io_outWtPS(PEs_3_7_io_outWtPS),
    .io_outAct(PEs_3_7_io_outAct),
    .io_inwtValid(PEs_3_7_io_inwtValid)
  );
  PE PEs_4_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_0_clock),
    .io_inAct(PEs_4_0_io_inAct),
    .io_inWtPS(PEs_4_0_io_inWtPS),
    .io_outWtPS(PEs_4_0_io_outWtPS),
    .io_outAct(PEs_4_0_io_outAct),
    .io_inwtValid(PEs_4_0_io_inwtValid)
  );
  PE PEs_4_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_1_clock),
    .io_inAct(PEs_4_1_io_inAct),
    .io_inWtPS(PEs_4_1_io_inWtPS),
    .io_outWtPS(PEs_4_1_io_outWtPS),
    .io_outAct(PEs_4_1_io_outAct),
    .io_inwtValid(PEs_4_1_io_inwtValid)
  );
  PE PEs_4_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_2_clock),
    .io_inAct(PEs_4_2_io_inAct),
    .io_inWtPS(PEs_4_2_io_inWtPS),
    .io_outWtPS(PEs_4_2_io_outWtPS),
    .io_outAct(PEs_4_2_io_outAct),
    .io_inwtValid(PEs_4_2_io_inwtValid)
  );
  PE PEs_4_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_3_clock),
    .io_inAct(PEs_4_3_io_inAct),
    .io_inWtPS(PEs_4_3_io_inWtPS),
    .io_outWtPS(PEs_4_3_io_outWtPS),
    .io_outAct(PEs_4_3_io_outAct),
    .io_inwtValid(PEs_4_3_io_inwtValid)
  );
  PE PEs_4_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_4_clock),
    .io_inAct(PEs_4_4_io_inAct),
    .io_inWtPS(PEs_4_4_io_inWtPS),
    .io_outWtPS(PEs_4_4_io_outWtPS),
    .io_outAct(PEs_4_4_io_outAct),
    .io_inwtValid(PEs_4_4_io_inwtValid)
  );
  PE PEs_4_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_5_clock),
    .io_inAct(PEs_4_5_io_inAct),
    .io_inWtPS(PEs_4_5_io_inWtPS),
    .io_outWtPS(PEs_4_5_io_outWtPS),
    .io_outAct(PEs_4_5_io_outAct),
    .io_inwtValid(PEs_4_5_io_inwtValid)
  );
  PE PEs_4_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_6_clock),
    .io_inAct(PEs_4_6_io_inAct),
    .io_inWtPS(PEs_4_6_io_inWtPS),
    .io_outWtPS(PEs_4_6_io_outWtPS),
    .io_outAct(PEs_4_6_io_outAct),
    .io_inwtValid(PEs_4_6_io_inwtValid)
  );
  PE PEs_4_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_4_7_clock),
    .io_inAct(PEs_4_7_io_inAct),
    .io_inWtPS(PEs_4_7_io_inWtPS),
    .io_outWtPS(PEs_4_7_io_outWtPS),
    .io_outAct(PEs_4_7_io_outAct),
    .io_inwtValid(PEs_4_7_io_inwtValid)
  );
  PE PEs_5_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_0_clock),
    .io_inAct(PEs_5_0_io_inAct),
    .io_inWtPS(PEs_5_0_io_inWtPS),
    .io_outWtPS(PEs_5_0_io_outWtPS),
    .io_outAct(PEs_5_0_io_outAct),
    .io_inwtValid(PEs_5_0_io_inwtValid)
  );
  PE PEs_5_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_1_clock),
    .io_inAct(PEs_5_1_io_inAct),
    .io_inWtPS(PEs_5_1_io_inWtPS),
    .io_outWtPS(PEs_5_1_io_outWtPS),
    .io_outAct(PEs_5_1_io_outAct),
    .io_inwtValid(PEs_5_1_io_inwtValid)
  );
  PE PEs_5_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_2_clock),
    .io_inAct(PEs_5_2_io_inAct),
    .io_inWtPS(PEs_5_2_io_inWtPS),
    .io_outWtPS(PEs_5_2_io_outWtPS),
    .io_outAct(PEs_5_2_io_outAct),
    .io_inwtValid(PEs_5_2_io_inwtValid)
  );
  PE PEs_5_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_3_clock),
    .io_inAct(PEs_5_3_io_inAct),
    .io_inWtPS(PEs_5_3_io_inWtPS),
    .io_outWtPS(PEs_5_3_io_outWtPS),
    .io_outAct(PEs_5_3_io_outAct),
    .io_inwtValid(PEs_5_3_io_inwtValid)
  );
  PE PEs_5_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_4_clock),
    .io_inAct(PEs_5_4_io_inAct),
    .io_inWtPS(PEs_5_4_io_inWtPS),
    .io_outWtPS(PEs_5_4_io_outWtPS),
    .io_outAct(PEs_5_4_io_outAct),
    .io_inwtValid(PEs_5_4_io_inwtValid)
  );
  PE PEs_5_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_5_clock),
    .io_inAct(PEs_5_5_io_inAct),
    .io_inWtPS(PEs_5_5_io_inWtPS),
    .io_outWtPS(PEs_5_5_io_outWtPS),
    .io_outAct(PEs_5_5_io_outAct),
    .io_inwtValid(PEs_5_5_io_inwtValid)
  );
  PE PEs_5_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_6_clock),
    .io_inAct(PEs_5_6_io_inAct),
    .io_inWtPS(PEs_5_6_io_inWtPS),
    .io_outWtPS(PEs_5_6_io_outWtPS),
    .io_outAct(PEs_5_6_io_outAct),
    .io_inwtValid(PEs_5_6_io_inwtValid)
  );
  PE PEs_5_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_5_7_clock),
    .io_inAct(PEs_5_7_io_inAct),
    .io_inWtPS(PEs_5_7_io_inWtPS),
    .io_outWtPS(PEs_5_7_io_outWtPS),
    .io_outAct(PEs_5_7_io_outAct),
    .io_inwtValid(PEs_5_7_io_inwtValid)
  );
  PE PEs_6_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_0_clock),
    .io_inAct(PEs_6_0_io_inAct),
    .io_inWtPS(PEs_6_0_io_inWtPS),
    .io_outWtPS(PEs_6_0_io_outWtPS),
    .io_outAct(PEs_6_0_io_outAct),
    .io_inwtValid(PEs_6_0_io_inwtValid)
  );
  PE PEs_6_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_1_clock),
    .io_inAct(PEs_6_1_io_inAct),
    .io_inWtPS(PEs_6_1_io_inWtPS),
    .io_outWtPS(PEs_6_1_io_outWtPS),
    .io_outAct(PEs_6_1_io_outAct),
    .io_inwtValid(PEs_6_1_io_inwtValid)
  );
  PE PEs_6_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_2_clock),
    .io_inAct(PEs_6_2_io_inAct),
    .io_inWtPS(PEs_6_2_io_inWtPS),
    .io_outWtPS(PEs_6_2_io_outWtPS),
    .io_outAct(PEs_6_2_io_outAct),
    .io_inwtValid(PEs_6_2_io_inwtValid)
  );
  PE PEs_6_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_3_clock),
    .io_inAct(PEs_6_3_io_inAct),
    .io_inWtPS(PEs_6_3_io_inWtPS),
    .io_outWtPS(PEs_6_3_io_outWtPS),
    .io_outAct(PEs_6_3_io_outAct),
    .io_inwtValid(PEs_6_3_io_inwtValid)
  );
  PE PEs_6_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_4_clock),
    .io_inAct(PEs_6_4_io_inAct),
    .io_inWtPS(PEs_6_4_io_inWtPS),
    .io_outWtPS(PEs_6_4_io_outWtPS),
    .io_outAct(PEs_6_4_io_outAct),
    .io_inwtValid(PEs_6_4_io_inwtValid)
  );
  PE PEs_6_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_5_clock),
    .io_inAct(PEs_6_5_io_inAct),
    .io_inWtPS(PEs_6_5_io_inWtPS),
    .io_outWtPS(PEs_6_5_io_outWtPS),
    .io_outAct(PEs_6_5_io_outAct),
    .io_inwtValid(PEs_6_5_io_inwtValid)
  );
  PE PEs_6_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_6_clock),
    .io_inAct(PEs_6_6_io_inAct),
    .io_inWtPS(PEs_6_6_io_inWtPS),
    .io_outWtPS(PEs_6_6_io_outWtPS),
    .io_outAct(PEs_6_6_io_outAct),
    .io_inwtValid(PEs_6_6_io_inwtValid)
  );
  PE PEs_6_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_6_7_clock),
    .io_inAct(PEs_6_7_io_inAct),
    .io_inWtPS(PEs_6_7_io_inWtPS),
    .io_outWtPS(PEs_6_7_io_outWtPS),
    .io_outAct(PEs_6_7_io_outAct),
    .io_inwtValid(PEs_6_7_io_inwtValid)
  );
  PE PEs_7_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_0_clock),
    .io_inAct(PEs_7_0_io_inAct),
    .io_inWtPS(PEs_7_0_io_inWtPS),
    .io_outWtPS(PEs_7_0_io_outWtPS),
    .io_outAct(PEs_7_0_io_outAct),
    .io_inwtValid(PEs_7_0_io_inwtValid)
  );
  PE PEs_7_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_1_clock),
    .io_inAct(PEs_7_1_io_inAct),
    .io_inWtPS(PEs_7_1_io_inWtPS),
    .io_outWtPS(PEs_7_1_io_outWtPS),
    .io_outAct(PEs_7_1_io_outAct),
    .io_inwtValid(PEs_7_1_io_inwtValid)
  );
  PE PEs_7_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_2_clock),
    .io_inAct(PEs_7_2_io_inAct),
    .io_inWtPS(PEs_7_2_io_inWtPS),
    .io_outWtPS(PEs_7_2_io_outWtPS),
    .io_outAct(PEs_7_2_io_outAct),
    .io_inwtValid(PEs_7_2_io_inwtValid)
  );
  PE PEs_7_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_3_clock),
    .io_inAct(PEs_7_3_io_inAct),
    .io_inWtPS(PEs_7_3_io_inWtPS),
    .io_outWtPS(PEs_7_3_io_outWtPS),
    .io_outAct(PEs_7_3_io_outAct),
    .io_inwtValid(PEs_7_3_io_inwtValid)
  );
  PE PEs_7_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_4_clock),
    .io_inAct(PEs_7_4_io_inAct),
    .io_inWtPS(PEs_7_4_io_inWtPS),
    .io_outWtPS(PEs_7_4_io_outWtPS),
    .io_outAct(PEs_7_4_io_outAct),
    .io_inwtValid(PEs_7_4_io_inwtValid)
  );
  PE PEs_7_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_5_clock),
    .io_inAct(PEs_7_5_io_inAct),
    .io_inWtPS(PEs_7_5_io_inWtPS),
    .io_outWtPS(PEs_7_5_io_outWtPS),
    .io_outAct(PEs_7_5_io_outAct),
    .io_inwtValid(PEs_7_5_io_inwtValid)
  );
  PE PEs_7_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_6_clock),
    .io_inAct(PEs_7_6_io_inAct),
    .io_inWtPS(PEs_7_6_io_inWtPS),
    .io_outWtPS(PEs_7_6_io_outWtPS),
    .io_outAct(PEs_7_6_io_outAct),
    .io_inwtValid(PEs_7_6_io_inwtValid)
  );
  PE PEs_7_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_7_7_clock),
    .io_inAct(PEs_7_7_io_inAct),
    .io_inWtPS(PEs_7_7_io_inWtPS),
    .io_outWtPS(PEs_7_7_io_outWtPS),
    .io_outAct(PEs_7_7_io_outAct),
    .io_inwtValid(PEs_7_7_io_inwtValid)
  );
  PE PEs_8_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_0_clock),
    .io_inAct(PEs_8_0_io_inAct),
    .io_inWtPS(PEs_8_0_io_inWtPS),
    .io_outWtPS(PEs_8_0_io_outWtPS),
    .io_outAct(PEs_8_0_io_outAct),
    .io_inwtValid(PEs_8_0_io_inwtValid)
  );
  PE PEs_8_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_1_clock),
    .io_inAct(PEs_8_1_io_inAct),
    .io_inWtPS(PEs_8_1_io_inWtPS),
    .io_outWtPS(PEs_8_1_io_outWtPS),
    .io_outAct(PEs_8_1_io_outAct),
    .io_inwtValid(PEs_8_1_io_inwtValid)
  );
  PE PEs_8_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_2_clock),
    .io_inAct(PEs_8_2_io_inAct),
    .io_inWtPS(PEs_8_2_io_inWtPS),
    .io_outWtPS(PEs_8_2_io_outWtPS),
    .io_outAct(PEs_8_2_io_outAct),
    .io_inwtValid(PEs_8_2_io_inwtValid)
  );
  PE PEs_8_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_3_clock),
    .io_inAct(PEs_8_3_io_inAct),
    .io_inWtPS(PEs_8_3_io_inWtPS),
    .io_outWtPS(PEs_8_3_io_outWtPS),
    .io_outAct(PEs_8_3_io_outAct),
    .io_inwtValid(PEs_8_3_io_inwtValid)
  );
  PE PEs_8_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_4_clock),
    .io_inAct(PEs_8_4_io_inAct),
    .io_inWtPS(PEs_8_4_io_inWtPS),
    .io_outWtPS(PEs_8_4_io_outWtPS),
    .io_outAct(PEs_8_4_io_outAct),
    .io_inwtValid(PEs_8_4_io_inwtValid)
  );
  PE PEs_8_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_5_clock),
    .io_inAct(PEs_8_5_io_inAct),
    .io_inWtPS(PEs_8_5_io_inWtPS),
    .io_outWtPS(PEs_8_5_io_outWtPS),
    .io_outAct(PEs_8_5_io_outAct),
    .io_inwtValid(PEs_8_5_io_inwtValid)
  );
  PE PEs_8_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_6_clock),
    .io_inAct(PEs_8_6_io_inAct),
    .io_inWtPS(PEs_8_6_io_inWtPS),
    .io_outWtPS(PEs_8_6_io_outWtPS),
    .io_outAct(PEs_8_6_io_outAct),
    .io_inwtValid(PEs_8_6_io_inwtValid)
  );
  PE PEs_8_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_8_7_clock),
    .io_inAct(PEs_8_7_io_inAct),
    .io_inWtPS(PEs_8_7_io_inWtPS),
    .io_outWtPS(PEs_8_7_io_outWtPS),
    .io_outAct(PEs_8_7_io_outAct),
    .io_inwtValid(PEs_8_7_io_inwtValid)
  );
  PE PEs_9_0 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_0_clock),
    .io_inAct(PEs_9_0_io_inAct),
    .io_inWtPS(PEs_9_0_io_inWtPS),
    .io_outWtPS(PEs_9_0_io_outWtPS),
    .io_outAct(PEs_9_0_io_outAct),
    .io_inwtValid(PEs_9_0_io_inwtValid)
  );
  PE PEs_9_1 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_1_clock),
    .io_inAct(PEs_9_1_io_inAct),
    .io_inWtPS(PEs_9_1_io_inWtPS),
    .io_outWtPS(PEs_9_1_io_outWtPS),
    .io_outAct(PEs_9_1_io_outAct),
    .io_inwtValid(PEs_9_1_io_inwtValid)
  );
  PE PEs_9_2 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_2_clock),
    .io_inAct(PEs_9_2_io_inAct),
    .io_inWtPS(PEs_9_2_io_inWtPS),
    .io_outWtPS(PEs_9_2_io_outWtPS),
    .io_outAct(PEs_9_2_io_outAct),
    .io_inwtValid(PEs_9_2_io_inwtValid)
  );
  PE PEs_9_3 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_3_clock),
    .io_inAct(PEs_9_3_io_inAct),
    .io_inWtPS(PEs_9_3_io_inWtPS),
    .io_outWtPS(PEs_9_3_io_outWtPS),
    .io_outAct(PEs_9_3_io_outAct),
    .io_inwtValid(PEs_9_3_io_inwtValid)
  );
  PE PEs_9_4 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_4_clock),
    .io_inAct(PEs_9_4_io_inAct),
    .io_inWtPS(PEs_9_4_io_inWtPS),
    .io_outWtPS(PEs_9_4_io_outWtPS),
    .io_outAct(PEs_9_4_io_outAct),
    .io_inwtValid(PEs_9_4_io_inwtValid)
  );
  PE PEs_9_5 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_5_clock),
    .io_inAct(PEs_9_5_io_inAct),
    .io_inWtPS(PEs_9_5_io_inWtPS),
    .io_outWtPS(PEs_9_5_io_outWtPS),
    .io_outAct(PEs_9_5_io_outAct),
    .io_inwtValid(PEs_9_5_io_inwtValid)
  );
  PE PEs_9_6 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_6_clock),
    .io_inAct(PEs_9_6_io_inAct),
    .io_inWtPS(PEs_9_6_io_inWtPS),
    .io_outWtPS(PEs_9_6_io_outWtPS),
    .io_outAct(PEs_9_6_io_outAct),
    .io_inwtValid(PEs_9_6_io_inwtValid)
  );
  PE PEs_9_7 ( // @[SystolicArray.scala 18:65]
    .clock(PEs_9_7_clock),
    .io_inAct(PEs_9_7_io_inAct),
    .io_inWtPS(PEs_9_7_io_inWtPS),
    .io_outWtPS(PEs_9_7_io_outWtPS),
    .io_outAct(PEs_9_7_io_outAct),
    .io_inwtValid(PEs_9_7_io_inwtValid)
  );
  assign io_outSum_0 = PEs_9_0_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_1 = PEs_9_1_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_2 = PEs_9_2_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_3 = PEs_9_3_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_4 = PEs_9_4_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_5 = PEs_9_5_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_6 = PEs_9_6_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign io_outSum_7 = PEs_9_7_io_outWtPS; // @[SystolicArray.scala 35:46]
  assign PEs_0_0_clock = clock;
  assign PEs_0_0_io_inAct = io_inAct_0; // @[SystolicArray.scala 38:44]
  assign PEs_0_0_io_inWtPS = {{24{io_inWeight_0[15]}},io_inWeight_0}; // @[SystolicArray.scala 31:45]
  assign PEs_0_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_1_clock = clock;
  assign PEs_0_1_io_inAct = PEs_0_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_1_io_inWtPS = {{24{io_inWeight_1[15]}},io_inWeight_1}; // @[SystolicArray.scala 31:45]
  assign PEs_0_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_2_clock = clock;
  assign PEs_0_2_io_inAct = PEs_0_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_2_io_inWtPS = {{24{io_inWeight_2[15]}},io_inWeight_2}; // @[SystolicArray.scala 31:45]
  assign PEs_0_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_3_clock = clock;
  assign PEs_0_3_io_inAct = PEs_0_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_3_io_inWtPS = {{24{io_inWeight_3[15]}},io_inWeight_3}; // @[SystolicArray.scala 31:45]
  assign PEs_0_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_4_clock = clock;
  assign PEs_0_4_io_inAct = PEs_0_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_4_io_inWtPS = {{24{io_inWeight_4[15]}},io_inWeight_4}; // @[SystolicArray.scala 31:45]
  assign PEs_0_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_5_clock = clock;
  assign PEs_0_5_io_inAct = PEs_0_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_5_io_inWtPS = {{24{io_inWeight_5[15]}},io_inWeight_5}; // @[SystolicArray.scala 31:45]
  assign PEs_0_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_6_clock = clock;
  assign PEs_0_6_io_inAct = PEs_0_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_6_io_inWtPS = {{24{io_inWeight_6[15]}},io_inWeight_6}; // @[SystolicArray.scala 31:45]
  assign PEs_0_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_0_7_clock = clock;
  assign PEs_0_7_io_inAct = PEs_0_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_0_7_io_inWtPS = {{24{io_inWeight_7[15]}},io_inWeight_7}; // @[SystolicArray.scala 31:45]
  assign PEs_0_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_0_clock = clock;
  assign PEs_1_0_io_inAct = io_inAct_1; // @[SystolicArray.scala 38:44]
  assign PEs_1_0_io_inWtPS = PEs_0_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_1_clock = clock;
  assign PEs_1_1_io_inAct = PEs_1_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_1_io_inWtPS = PEs_0_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_2_clock = clock;
  assign PEs_1_2_io_inAct = PEs_1_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_2_io_inWtPS = PEs_0_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_3_clock = clock;
  assign PEs_1_3_io_inAct = PEs_1_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_3_io_inWtPS = PEs_0_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_4_clock = clock;
  assign PEs_1_4_io_inAct = PEs_1_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_4_io_inWtPS = PEs_0_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_5_clock = clock;
  assign PEs_1_5_io_inAct = PEs_1_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_5_io_inWtPS = PEs_0_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_6_clock = clock;
  assign PEs_1_6_io_inAct = PEs_1_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_6_io_inWtPS = PEs_0_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_1_7_clock = clock;
  assign PEs_1_7_io_inAct = PEs_1_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_1_7_io_inWtPS = PEs_0_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_1_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_0_clock = clock;
  assign PEs_2_0_io_inAct = io_inAct_2; // @[SystolicArray.scala 38:44]
  assign PEs_2_0_io_inWtPS = PEs_1_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_1_clock = clock;
  assign PEs_2_1_io_inAct = PEs_2_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_1_io_inWtPS = PEs_1_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_2_clock = clock;
  assign PEs_2_2_io_inAct = PEs_2_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_2_io_inWtPS = PEs_1_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_3_clock = clock;
  assign PEs_2_3_io_inAct = PEs_2_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_3_io_inWtPS = PEs_1_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_4_clock = clock;
  assign PEs_2_4_io_inAct = PEs_2_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_4_io_inWtPS = PEs_1_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_5_clock = clock;
  assign PEs_2_5_io_inAct = PEs_2_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_5_io_inWtPS = PEs_1_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_6_clock = clock;
  assign PEs_2_6_io_inAct = PEs_2_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_6_io_inWtPS = PEs_1_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_2_7_clock = clock;
  assign PEs_2_7_io_inAct = PEs_2_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_2_7_io_inWtPS = PEs_1_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_2_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_0_clock = clock;
  assign PEs_3_0_io_inAct = io_inAct_3; // @[SystolicArray.scala 38:44]
  assign PEs_3_0_io_inWtPS = PEs_2_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_1_clock = clock;
  assign PEs_3_1_io_inAct = PEs_3_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_1_io_inWtPS = PEs_2_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_2_clock = clock;
  assign PEs_3_2_io_inAct = PEs_3_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_2_io_inWtPS = PEs_2_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_3_clock = clock;
  assign PEs_3_3_io_inAct = PEs_3_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_3_io_inWtPS = PEs_2_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_4_clock = clock;
  assign PEs_3_4_io_inAct = PEs_3_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_4_io_inWtPS = PEs_2_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_5_clock = clock;
  assign PEs_3_5_io_inAct = PEs_3_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_5_io_inWtPS = PEs_2_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_6_clock = clock;
  assign PEs_3_6_io_inAct = PEs_3_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_6_io_inWtPS = PEs_2_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_3_7_clock = clock;
  assign PEs_3_7_io_inAct = PEs_3_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_3_7_io_inWtPS = PEs_2_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_3_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_0_clock = clock;
  assign PEs_4_0_io_inAct = io_inAct_4; // @[SystolicArray.scala 38:44]
  assign PEs_4_0_io_inWtPS = PEs_3_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_1_clock = clock;
  assign PEs_4_1_io_inAct = PEs_4_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_1_io_inWtPS = PEs_3_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_2_clock = clock;
  assign PEs_4_2_io_inAct = PEs_4_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_2_io_inWtPS = PEs_3_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_3_clock = clock;
  assign PEs_4_3_io_inAct = PEs_4_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_3_io_inWtPS = PEs_3_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_4_clock = clock;
  assign PEs_4_4_io_inAct = PEs_4_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_4_io_inWtPS = PEs_3_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_5_clock = clock;
  assign PEs_4_5_io_inAct = PEs_4_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_5_io_inWtPS = PEs_3_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_6_clock = clock;
  assign PEs_4_6_io_inAct = PEs_4_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_6_io_inWtPS = PEs_3_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_4_7_clock = clock;
  assign PEs_4_7_io_inAct = PEs_4_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_4_7_io_inWtPS = PEs_3_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_4_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_0_clock = clock;
  assign PEs_5_0_io_inAct = io_inAct_5; // @[SystolicArray.scala 38:44]
  assign PEs_5_0_io_inWtPS = PEs_4_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_1_clock = clock;
  assign PEs_5_1_io_inAct = PEs_5_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_1_io_inWtPS = PEs_4_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_2_clock = clock;
  assign PEs_5_2_io_inAct = PEs_5_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_2_io_inWtPS = PEs_4_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_3_clock = clock;
  assign PEs_5_3_io_inAct = PEs_5_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_3_io_inWtPS = PEs_4_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_4_clock = clock;
  assign PEs_5_4_io_inAct = PEs_5_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_4_io_inWtPS = PEs_4_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_5_clock = clock;
  assign PEs_5_5_io_inAct = PEs_5_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_5_io_inWtPS = PEs_4_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_6_clock = clock;
  assign PEs_5_6_io_inAct = PEs_5_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_6_io_inWtPS = PEs_4_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_5_7_clock = clock;
  assign PEs_5_7_io_inAct = PEs_5_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_5_7_io_inWtPS = PEs_4_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_5_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_0_clock = clock;
  assign PEs_6_0_io_inAct = io_inAct_6; // @[SystolicArray.scala 38:44]
  assign PEs_6_0_io_inWtPS = PEs_5_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_1_clock = clock;
  assign PEs_6_1_io_inAct = PEs_6_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_1_io_inWtPS = PEs_5_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_2_clock = clock;
  assign PEs_6_2_io_inAct = PEs_6_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_2_io_inWtPS = PEs_5_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_3_clock = clock;
  assign PEs_6_3_io_inAct = PEs_6_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_3_io_inWtPS = PEs_5_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_4_clock = clock;
  assign PEs_6_4_io_inAct = PEs_6_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_4_io_inWtPS = PEs_5_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_5_clock = clock;
  assign PEs_6_5_io_inAct = PEs_6_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_5_io_inWtPS = PEs_5_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_6_clock = clock;
  assign PEs_6_6_io_inAct = PEs_6_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_6_io_inWtPS = PEs_5_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_6_7_clock = clock;
  assign PEs_6_7_io_inAct = PEs_6_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_6_7_io_inWtPS = PEs_5_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_6_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_0_clock = clock;
  assign PEs_7_0_io_inAct = io_inAct_7; // @[SystolicArray.scala 38:44]
  assign PEs_7_0_io_inWtPS = PEs_6_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_1_clock = clock;
  assign PEs_7_1_io_inAct = PEs_7_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_1_io_inWtPS = PEs_6_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_2_clock = clock;
  assign PEs_7_2_io_inAct = PEs_7_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_2_io_inWtPS = PEs_6_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_3_clock = clock;
  assign PEs_7_3_io_inAct = PEs_7_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_3_io_inWtPS = PEs_6_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_4_clock = clock;
  assign PEs_7_4_io_inAct = PEs_7_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_4_io_inWtPS = PEs_6_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_5_clock = clock;
  assign PEs_7_5_io_inAct = PEs_7_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_5_io_inWtPS = PEs_6_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_6_clock = clock;
  assign PEs_7_6_io_inAct = PEs_7_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_6_io_inWtPS = PEs_6_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_7_7_clock = clock;
  assign PEs_7_7_io_inAct = PEs_7_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_7_7_io_inWtPS = PEs_6_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_7_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_0_clock = clock;
  assign PEs_8_0_io_inAct = io_inAct_8; // @[SystolicArray.scala 38:44]
  assign PEs_8_0_io_inWtPS = PEs_7_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_1_clock = clock;
  assign PEs_8_1_io_inAct = PEs_8_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_1_io_inWtPS = PEs_7_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_2_clock = clock;
  assign PEs_8_2_io_inAct = PEs_8_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_2_io_inWtPS = PEs_7_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_3_clock = clock;
  assign PEs_8_3_io_inAct = PEs_8_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_3_io_inWtPS = PEs_7_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_4_clock = clock;
  assign PEs_8_4_io_inAct = PEs_8_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_4_io_inWtPS = PEs_7_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_5_clock = clock;
  assign PEs_8_5_io_inAct = PEs_8_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_5_io_inWtPS = PEs_7_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_6_clock = clock;
  assign PEs_8_6_io_inAct = PEs_8_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_6_io_inWtPS = PEs_7_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_8_7_clock = clock;
  assign PEs_8_7_io_inAct = PEs_8_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_8_7_io_inWtPS = PEs_7_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_8_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_0_clock = clock;
  assign PEs_9_0_io_inAct = io_inAct_9; // @[SystolicArray.scala 38:44]
  assign PEs_9_0_io_inWtPS = PEs_8_0_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_0_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_1_clock = clock;
  assign PEs_9_1_io_inAct = PEs_9_0_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_1_io_inWtPS = PEs_8_1_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_1_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_2_clock = clock;
  assign PEs_9_2_io_inAct = PEs_9_1_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_2_io_inWtPS = PEs_8_2_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_2_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_3_clock = clock;
  assign PEs_9_3_io_inAct = PEs_9_2_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_3_io_inWtPS = PEs_8_3_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_3_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_4_clock = clock;
  assign PEs_9_4_io_inAct = PEs_9_3_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_4_io_inWtPS = PEs_8_4_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_4_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_5_clock = clock;
  assign PEs_9_5_io_inAct = PEs_9_4_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_5_io_inWtPS = PEs_8_5_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_5_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_6_clock = clock;
  assign PEs_9_6_io_inAct = PEs_9_5_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_6_io_inWtPS = PEs_8_6_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_6_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  assign PEs_9_7_clock = clock;
  assign PEs_9_7_io_inAct = PEs_9_6_io_outAct; // @[SystolicArray.scala 39:44]
  assign PEs_9_7_io_inWtPS = PEs_8_7_io_outWtPS; // @[SystolicArray.scala 32:45]
  assign PEs_9_7_io_inwtValid = validReg; // @[SystolicArray.scala 25:40]
  always @(posedge clock) begin
    validReg <= io_inwtValid; // @[SystolicArray.scala 22:25]
  end
endmodule
module BiasActivation(
  input         clock,
  input  [39:0] io_inSum_0,
  input  [39:0] io_inSum_1,
  input  [39:0] io_inSum_2,
  input  [39:0] io_inSum_3,
  input  [39:0] io_inSum_4,
  input  [39:0] io_inSum_5,
  input  [39:0] io_inSum_6,
  input  [39:0] io_inSum_7,
  input  [39:0] io_inSum_8,
  input  [39:0] io_inSum_9,
  output [15:0] io_outAct_0,
  output [15:0] io_outAct_1,
  output [15:0] io_outAct_2,
  output [15:0] io_outAct_3,
  output [15:0] io_outAct_4,
  output [15:0] io_outAct_5,
  output [15:0] io_outAct_6,
  output [15:0] io_outAct_7,
  output [15:0] io_outAct_8,
  output [15:0] io_outAct_9,
  input  [15:0] io_inBias_0,
  input  [15:0] io_inBias_1,
  input  [15:0] io_inBias_2,
  input  [15:0] io_inBias_3,
  input  [15:0] io_inBias_4,
  input  [15:0] io_inBias_5,
  input  [15:0] io_inBias_6,
  input  [15:0] io_inBias_7,
  input  [15:0] io_inBias_8,
  input  [15:0] io_inBias_9,
  input         io_inBiasValid
);
  reg [15:0] biasReg_0; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_1; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_2; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_3; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_4; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_5; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_6; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_7; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_8; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_9; // @[BiasActivation.scala 28:22]
  reg [39:0] plusReg_0; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_1; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_2; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_3; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_4; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_5; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_6; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_7; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_8; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_9; // @[BiasActivation.scala 29:22]
  reg [15:0] actReg_0; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_1; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_2; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_3; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_4; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_5; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_6; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_7; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_8; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_9; // @[BiasActivation.scala 30:22]
  reg  sumReg_0; // @[BiasActivation.scala 31:22]
  reg  sumReg_1; // @[BiasActivation.scala 31:22]
  reg  sumReg_2; // @[BiasActivation.scala 31:22]
  reg  sumReg_3; // @[BiasActivation.scala 31:22]
  reg  sumReg_4; // @[BiasActivation.scala 31:22]
  reg  sumReg_5; // @[BiasActivation.scala 31:22]
  reg  sumReg_6; // @[BiasActivation.scala 31:22]
  reg  sumReg_7; // @[BiasActivation.scala 31:22]
  reg  sumReg_8; // @[BiasActivation.scala 31:22]
  reg  sumReg_9; // @[BiasActivation.scala 31:22]
  reg  validReg; // @[BiasActivation.scala 32:26]
  wire [29:0] _T = {$signed(biasReg_0), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_30 = {{10{_T[29]}},_T}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_4 = {$signed(biasReg_1), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_31 = {{10{_T_4[29]}},_T_4}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_8 = {$signed(biasReg_2), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_32 = {{10{_T_8[29]}},_T_8}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_12 = {$signed(biasReg_3), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_33 = {{10{_T_12[29]}},_T_12}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_16 = {$signed(biasReg_4), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_34 = {{10{_T_16[29]}},_T_16}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_20 = {$signed(biasReg_5), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_35 = {{10{_T_20[29]}},_T_20}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_24 = {$signed(biasReg_6), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_36 = {{10{_T_24[29]}},_T_24}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_28 = {$signed(biasReg_7), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_37 = {{10{_T_28[29]}},_T_28}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_32 = {$signed(biasReg_8), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_38 = {{10{_T_32[29]}},_T_32}; // @[BiasActivation.scala 56:80]
  wire [29:0] _T_36 = {$signed(biasReg_9), 14'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_39 = {{10{_T_36[29]}},_T_36}; // @[BiasActivation.scala 56:80]
  wire [15:0] _truncWire_0_T_1 = plusReg_0[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_10 = plusReg_0[30] & ~sumReg_0 & ~biasReg_0[15] ? $signed(16'sh8000) : $signed(_truncWire_0_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_0 = ~plusReg_0[30] & sumReg_0 & biasReg_0[15] ? $signed(16'sh7fff) : $signed(_GEN_10); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_1_T_1 = plusReg_1[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_12 = plusReg_1[30] & ~sumReg_1 & ~biasReg_1[15] ? $signed(16'sh8000) : $signed(_truncWire_1_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_1 = ~plusReg_1[30] & sumReg_1 & biasReg_1[15] ? $signed(16'sh7fff) : $signed(_GEN_12); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_2_T_1 = plusReg_2[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_14 = plusReg_2[30] & ~sumReg_2 & ~biasReg_2[15] ? $signed(16'sh8000) : $signed(_truncWire_2_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_2 = ~plusReg_2[30] & sumReg_2 & biasReg_2[15] ? $signed(16'sh7fff) : $signed(_GEN_14); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_3_T_1 = plusReg_3[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_16 = plusReg_3[30] & ~sumReg_3 & ~biasReg_3[15] ? $signed(16'sh8000) : $signed(_truncWire_3_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_3 = ~plusReg_3[30] & sumReg_3 & biasReg_3[15] ? $signed(16'sh7fff) : $signed(_GEN_16); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_4_T_1 = plusReg_4[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_18 = plusReg_4[30] & ~sumReg_4 & ~biasReg_4[15] ? $signed(16'sh8000) : $signed(_truncWire_4_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_4 = ~plusReg_4[30] & sumReg_4 & biasReg_4[15] ? $signed(16'sh7fff) : $signed(_GEN_18); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_5_T_1 = plusReg_5[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_20 = plusReg_5[30] & ~sumReg_5 & ~biasReg_5[15] ? $signed(16'sh8000) : $signed(_truncWire_5_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_5 = ~plusReg_5[30] & sumReg_5 & biasReg_5[15] ? $signed(16'sh7fff) : $signed(_GEN_20); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_6_T_1 = plusReg_6[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_22 = plusReg_6[30] & ~sumReg_6 & ~biasReg_6[15] ? $signed(16'sh8000) : $signed(_truncWire_6_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_6 = ~plusReg_6[30] & sumReg_6 & biasReg_6[15] ? $signed(16'sh7fff) : $signed(_GEN_22); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_7_T_1 = plusReg_7[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_24 = plusReg_7[30] & ~sumReg_7 & ~biasReg_7[15] ? $signed(16'sh8000) : $signed(_truncWire_7_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_7 = ~plusReg_7[30] & sumReg_7 & biasReg_7[15] ? $signed(16'sh7fff) : $signed(_GEN_24); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_8_T_1 = plusReg_8[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_26 = plusReg_8[30] & ~sumReg_8 & ~biasReg_8[15] ? $signed(16'sh8000) : $signed(_truncWire_8_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_8 = ~plusReg_8[30] & sumReg_8 & biasReg_8[15] ? $signed(16'sh7fff) : $signed(_GEN_26); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_9_T_1 = plusReg_9[30:15]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_28 = plusReg_9[30] & ~sumReg_9 & ~biasReg_9[15] ? $signed(16'sh8000) : $signed(_truncWire_9_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_9 = ~plusReg_9[30] & sumReg_9 & biasReg_9[15] ? $signed(16'sh7fff) : $signed(_GEN_28); // @[BiasActivation.scala 67:85 69:15]
  assign io_outAct_0 = actReg_0; // @[BiasActivation.scala 91:15]
  assign io_outAct_1 = actReg_1; // @[BiasActivation.scala 91:15]
  assign io_outAct_2 = actReg_2; // @[BiasActivation.scala 91:15]
  assign io_outAct_3 = actReg_3; // @[BiasActivation.scala 91:15]
  assign io_outAct_4 = actReg_4; // @[BiasActivation.scala 91:15]
  assign io_outAct_5 = actReg_5; // @[BiasActivation.scala 91:15]
  assign io_outAct_6 = actReg_6; // @[BiasActivation.scala 91:15]
  assign io_outAct_7 = actReg_7; // @[BiasActivation.scala 91:15]
  assign io_outAct_8 = actReg_8; // @[BiasActivation.scala 91:15]
  assign io_outAct_9 = actReg_9; // @[BiasActivation.scala 91:15]
  always @(posedge clock) begin
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_0 <= io_inBias_0; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_1 <= io_inBias_1; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_2 <= io_inBias_2; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_3 <= io_inBias_3; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_4 <= io_inBias_4; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_5 <= io_inBias_5; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_6 <= io_inBias_6; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_7 <= io_inBias_7; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_8 <= io_inBias_8; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_9 <= io_inBias_9; // @[BiasActivation.scala 50:17]
    end
    plusReg_0 <= $signed(_GEN_30) + $signed(io_inSum_0); // @[BiasActivation.scala 56:80]
    plusReg_1 <= $signed(_GEN_31) + $signed(io_inSum_1); // @[BiasActivation.scala 56:80]
    plusReg_2 <= $signed(_GEN_32) + $signed(io_inSum_2); // @[BiasActivation.scala 56:80]
    plusReg_3 <= $signed(_GEN_33) + $signed(io_inSum_3); // @[BiasActivation.scala 56:80]
    plusReg_4 <= $signed(_GEN_34) + $signed(io_inSum_4); // @[BiasActivation.scala 56:80]
    plusReg_5 <= $signed(_GEN_35) + $signed(io_inSum_5); // @[BiasActivation.scala 56:80]
    plusReg_6 <= $signed(_GEN_36) + $signed(io_inSum_6); // @[BiasActivation.scala 56:80]
    plusReg_7 <= $signed(_GEN_37) + $signed(io_inSum_7); // @[BiasActivation.scala 56:80]
    plusReg_8 <= $signed(_GEN_38) + $signed(io_inSum_8); // @[BiasActivation.scala 56:80]
    plusReg_9 <= $signed(_GEN_39) + $signed(io_inSum_9); // @[BiasActivation.scala 56:80]
    if ($signed(truncWire_0) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_0[30] & sumReg_0 & biasReg_0[15]) begin // @[BiasActivation.scala 67:85]
        actReg_0 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_0[30] & ~sumReg_0 & ~biasReg_0[15]) begin // @[BiasActivation.scala 70:92]
        actReg_0 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_0 <= _truncWire_0_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_0 <= 16'sh0;
    end
    if ($signed(truncWire_1) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_1[30] & sumReg_1 & biasReg_1[15]) begin // @[BiasActivation.scala 67:85]
        actReg_1 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_1[30] & ~sumReg_1 & ~biasReg_1[15]) begin // @[BiasActivation.scala 70:92]
        actReg_1 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_1 <= _truncWire_1_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_1 <= 16'sh0;
    end
    if ($signed(truncWire_2) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_2[30] & sumReg_2 & biasReg_2[15]) begin // @[BiasActivation.scala 67:85]
        actReg_2 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_2[30] & ~sumReg_2 & ~biasReg_2[15]) begin // @[BiasActivation.scala 70:92]
        actReg_2 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_2 <= _truncWire_2_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_2 <= 16'sh0;
    end
    if ($signed(truncWire_3) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_3[30] & sumReg_3 & biasReg_3[15]) begin // @[BiasActivation.scala 67:85]
        actReg_3 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_3[30] & ~sumReg_3 & ~biasReg_3[15]) begin // @[BiasActivation.scala 70:92]
        actReg_3 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_3 <= _truncWire_3_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_3 <= 16'sh0;
    end
    if ($signed(truncWire_4) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_4[30] & sumReg_4 & biasReg_4[15]) begin // @[BiasActivation.scala 67:85]
        actReg_4 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_4[30] & ~sumReg_4 & ~biasReg_4[15]) begin // @[BiasActivation.scala 70:92]
        actReg_4 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_4 <= _truncWire_4_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_4 <= 16'sh0;
    end
    if ($signed(truncWire_5) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_5[30] & sumReg_5 & biasReg_5[15]) begin // @[BiasActivation.scala 67:85]
        actReg_5 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_5[30] & ~sumReg_5 & ~biasReg_5[15]) begin // @[BiasActivation.scala 70:92]
        actReg_5 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_5 <= _truncWire_5_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_5 <= 16'sh0;
    end
    if ($signed(truncWire_6) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_6[30] & sumReg_6 & biasReg_6[15]) begin // @[BiasActivation.scala 67:85]
        actReg_6 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_6[30] & ~sumReg_6 & ~biasReg_6[15]) begin // @[BiasActivation.scala 70:92]
        actReg_6 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_6 <= _truncWire_6_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_6 <= 16'sh0;
    end
    if ($signed(truncWire_7) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_7[30] & sumReg_7 & biasReg_7[15]) begin // @[BiasActivation.scala 67:85]
        actReg_7 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_7[30] & ~sumReg_7 & ~biasReg_7[15]) begin // @[BiasActivation.scala 70:92]
        actReg_7 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_7 <= _truncWire_7_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_7 <= 16'sh0;
    end
    if ($signed(truncWire_8) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_8[30] & sumReg_8 & biasReg_8[15]) begin // @[BiasActivation.scala 67:85]
        actReg_8 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_8[30] & ~sumReg_8 & ~biasReg_8[15]) begin // @[BiasActivation.scala 70:92]
        actReg_8 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_8 <= _truncWire_8_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_8 <= 16'sh0;
    end
    if ($signed(truncWire_9) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_9[30] & sumReg_9 & biasReg_9[15]) begin // @[BiasActivation.scala 67:85]
        actReg_9 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_9[30] & ~sumReg_9 & ~biasReg_9[15]) begin // @[BiasActivation.scala 70:92]
        actReg_9 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_9 <= _truncWire_9_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_9 <= 16'sh0;
    end
    sumReg_0 <= io_inSum_0[30]; // @[BiasActivation.scala 61:59]
    sumReg_1 <= io_inSum_1[30]; // @[BiasActivation.scala 61:59]
    sumReg_2 <= io_inSum_2[30]; // @[BiasActivation.scala 61:59]
    sumReg_3 <= io_inSum_3[30]; // @[BiasActivation.scala 61:59]
    sumReg_4 <= io_inSum_4[30]; // @[BiasActivation.scala 61:59]
    sumReg_5 <= io_inSum_5[30]; // @[BiasActivation.scala 61:59]
    sumReg_6 <= io_inSum_6[30]; // @[BiasActivation.scala 61:59]
    sumReg_7 <= io_inSum_7[30]; // @[BiasActivation.scala 61:59]
    sumReg_8 <= io_inSum_8[30]; // @[BiasActivation.scala 61:59]
    sumReg_9 <= io_inSum_9[30]; // @[BiasActivation.scala 61:59]
    validReg <= io_inBiasValid; // @[BiasActivation.scala 32:26]
  end
endmodule
module BiasActivation_1(
  input         clock,
  input  [39:0] io_inSum_0,
  input  [39:0] io_inSum_1,
  input  [39:0] io_inSum_2,
  input  [39:0] io_inSum_3,
  input  [39:0] io_inSum_4,
  input  [39:0] io_inSum_5,
  input  [39:0] io_inSum_6,
  input  [39:0] io_inSum_7,
  input  [39:0] io_inSum_8,
  input  [39:0] io_inSum_9,
  output [15:0] io_outAct_0,
  output [15:0] io_outAct_1,
  output [15:0] io_outAct_2,
  output [15:0] io_outAct_3,
  output [15:0] io_outAct_4,
  output [15:0] io_outAct_5,
  output [15:0] io_outAct_6,
  output [15:0] io_outAct_7,
  output [15:0] io_outAct_8,
  output [15:0] io_outAct_9,
  input  [15:0] io_inBias_0,
  input  [15:0] io_inBias_1,
  input  [15:0] io_inBias_2,
  input  [15:0] io_inBias_3,
  input  [15:0] io_inBias_4,
  input  [15:0] io_inBias_5,
  input  [15:0] io_inBias_6,
  input  [15:0] io_inBias_7,
  input  [15:0] io_inBias_8,
  input  [15:0] io_inBias_9,
  input         io_inBiasValid
);
  reg [15:0] biasReg_0; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_1; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_2; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_3; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_4; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_5; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_6; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_7; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_8; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_9; // @[BiasActivation.scala 28:22]
  reg [39:0] plusReg_0; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_1; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_2; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_3; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_4; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_5; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_6; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_7; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_8; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_9; // @[BiasActivation.scala 29:22]
  reg [15:0] actReg_0; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_1; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_2; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_3; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_4; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_5; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_6; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_7; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_8; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_9; // @[BiasActivation.scala 30:22]
  reg  sumReg_0; // @[BiasActivation.scala 31:22]
  reg  sumReg_1; // @[BiasActivation.scala 31:22]
  reg  sumReg_2; // @[BiasActivation.scala 31:22]
  reg  sumReg_3; // @[BiasActivation.scala 31:22]
  reg  sumReg_4; // @[BiasActivation.scala 31:22]
  reg  sumReg_5; // @[BiasActivation.scala 31:22]
  reg  sumReg_6; // @[BiasActivation.scala 31:22]
  reg  sumReg_7; // @[BiasActivation.scala 31:22]
  reg  sumReg_8; // @[BiasActivation.scala 31:22]
  reg  sumReg_9; // @[BiasActivation.scala 31:22]
  reg  validReg; // @[BiasActivation.scala 32:26]
  wire [27:0] _T = {$signed(biasReg_0), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_30 = {{12{_T[27]}},_T}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_4 = {$signed(biasReg_1), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_31 = {{12{_T_4[27]}},_T_4}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_8 = {$signed(biasReg_2), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_32 = {{12{_T_8[27]}},_T_8}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_12 = {$signed(biasReg_3), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_33 = {{12{_T_12[27]}},_T_12}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_16 = {$signed(biasReg_4), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_34 = {{12{_T_16[27]}},_T_16}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_20 = {$signed(biasReg_5), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_35 = {{12{_T_20[27]}},_T_20}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_24 = {$signed(biasReg_6), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_36 = {{12{_T_24[27]}},_T_24}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_28 = {$signed(biasReg_7), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_37 = {{12{_T_28[27]}},_T_28}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_32 = {$signed(biasReg_8), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_38 = {{12{_T_32[27]}},_T_32}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_36 = {$signed(biasReg_9), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_39 = {{12{_T_36[27]}},_T_36}; // @[BiasActivation.scala 56:80]
  wire [15:0] _truncWire_0_T_1 = plusReg_0[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_10 = plusReg_0[28] & ~sumReg_0 & ~biasReg_0[15] ? $signed(16'sh8000) : $signed(_truncWire_0_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_0 = ~plusReg_0[28] & sumReg_0 & biasReg_0[15] ? $signed(16'sh7fff) : $signed(_GEN_10); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_1_T_1 = plusReg_1[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_12 = plusReg_1[28] & ~sumReg_1 & ~biasReg_1[15] ? $signed(16'sh8000) : $signed(_truncWire_1_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_1 = ~plusReg_1[28] & sumReg_1 & biasReg_1[15] ? $signed(16'sh7fff) : $signed(_GEN_12); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_2_T_1 = plusReg_2[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_14 = plusReg_2[28] & ~sumReg_2 & ~biasReg_2[15] ? $signed(16'sh8000) : $signed(_truncWire_2_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_2 = ~plusReg_2[28] & sumReg_2 & biasReg_2[15] ? $signed(16'sh7fff) : $signed(_GEN_14); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_3_T_1 = plusReg_3[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_16 = plusReg_3[28] & ~sumReg_3 & ~biasReg_3[15] ? $signed(16'sh8000) : $signed(_truncWire_3_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_3 = ~plusReg_3[28] & sumReg_3 & biasReg_3[15] ? $signed(16'sh7fff) : $signed(_GEN_16); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_4_T_1 = plusReg_4[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_18 = plusReg_4[28] & ~sumReg_4 & ~biasReg_4[15] ? $signed(16'sh8000) : $signed(_truncWire_4_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_4 = ~plusReg_4[28] & sumReg_4 & biasReg_4[15] ? $signed(16'sh7fff) : $signed(_GEN_18); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_5_T_1 = plusReg_5[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_20 = plusReg_5[28] & ~sumReg_5 & ~biasReg_5[15] ? $signed(16'sh8000) : $signed(_truncWire_5_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_5 = ~plusReg_5[28] & sumReg_5 & biasReg_5[15] ? $signed(16'sh7fff) : $signed(_GEN_20); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_6_T_1 = plusReg_6[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_22 = plusReg_6[28] & ~sumReg_6 & ~biasReg_6[15] ? $signed(16'sh8000) : $signed(_truncWire_6_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_6 = ~plusReg_6[28] & sumReg_6 & biasReg_6[15] ? $signed(16'sh7fff) : $signed(_GEN_22); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_7_T_1 = plusReg_7[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_24 = plusReg_7[28] & ~sumReg_7 & ~biasReg_7[15] ? $signed(16'sh8000) : $signed(_truncWire_7_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_7 = ~plusReg_7[28] & sumReg_7 & biasReg_7[15] ? $signed(16'sh7fff) : $signed(_GEN_24); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_8_T_1 = plusReg_8[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_26 = plusReg_8[28] & ~sumReg_8 & ~biasReg_8[15] ? $signed(16'sh8000) : $signed(_truncWire_8_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_8 = ~plusReg_8[28] & sumReg_8 & biasReg_8[15] ? $signed(16'sh7fff) : $signed(_GEN_26); // @[BiasActivation.scala 67:85 69:15]
  wire [15:0] _truncWire_9_T_1 = plusReg_9[28:13]; // @[BiasActivation.scala 74:66]
  wire [15:0] _GEN_28 = plusReg_9[28] & ~sumReg_9 & ~biasReg_9[15] ? $signed(16'sh8000) : $signed(_truncWire_9_T_1); // @[BiasActivation.scala 70:92 72:15 74:15]
  wire [15:0] truncWire_9 = ~plusReg_9[28] & sumReg_9 & biasReg_9[15] ? $signed(16'sh7fff) : $signed(_GEN_28); // @[BiasActivation.scala 67:85 69:15]
  assign io_outAct_0 = actReg_0; // @[BiasActivation.scala 91:15]
  assign io_outAct_1 = actReg_1; // @[BiasActivation.scala 91:15]
  assign io_outAct_2 = actReg_2; // @[BiasActivation.scala 91:15]
  assign io_outAct_3 = actReg_3; // @[BiasActivation.scala 91:15]
  assign io_outAct_4 = actReg_4; // @[BiasActivation.scala 91:15]
  assign io_outAct_5 = actReg_5; // @[BiasActivation.scala 91:15]
  assign io_outAct_6 = actReg_6; // @[BiasActivation.scala 91:15]
  assign io_outAct_7 = actReg_7; // @[BiasActivation.scala 91:15]
  assign io_outAct_8 = actReg_8; // @[BiasActivation.scala 91:15]
  assign io_outAct_9 = actReg_9; // @[BiasActivation.scala 91:15]
  always @(posedge clock) begin
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_0 <= io_inBias_0; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_1 <= io_inBias_1; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_2 <= io_inBias_2; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_3 <= io_inBias_3; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_4 <= io_inBias_4; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_5 <= io_inBias_5; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_6 <= io_inBias_6; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_7 <= io_inBias_7; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_8 <= io_inBias_8; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_9 <= io_inBias_9; // @[BiasActivation.scala 50:17]
    end
    plusReg_0 <= $signed(_GEN_30) + $signed(io_inSum_0); // @[BiasActivation.scala 56:80]
    plusReg_1 <= $signed(_GEN_31) + $signed(io_inSum_1); // @[BiasActivation.scala 56:80]
    plusReg_2 <= $signed(_GEN_32) + $signed(io_inSum_2); // @[BiasActivation.scala 56:80]
    plusReg_3 <= $signed(_GEN_33) + $signed(io_inSum_3); // @[BiasActivation.scala 56:80]
    plusReg_4 <= $signed(_GEN_34) + $signed(io_inSum_4); // @[BiasActivation.scala 56:80]
    plusReg_5 <= $signed(_GEN_35) + $signed(io_inSum_5); // @[BiasActivation.scala 56:80]
    plusReg_6 <= $signed(_GEN_36) + $signed(io_inSum_6); // @[BiasActivation.scala 56:80]
    plusReg_7 <= $signed(_GEN_37) + $signed(io_inSum_7); // @[BiasActivation.scala 56:80]
    plusReg_8 <= $signed(_GEN_38) + $signed(io_inSum_8); // @[BiasActivation.scala 56:80]
    plusReg_9 <= $signed(_GEN_39) + $signed(io_inSum_9); // @[BiasActivation.scala 56:80]
    if ($signed(truncWire_0) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_0[28] & sumReg_0 & biasReg_0[15]) begin // @[BiasActivation.scala 67:85]
        actReg_0 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_0[28] & ~sumReg_0 & ~biasReg_0[15]) begin // @[BiasActivation.scala 70:92]
        actReg_0 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_0 <= _truncWire_0_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_0 <= 16'sh0;
    end
    if ($signed(truncWire_1) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_1[28] & sumReg_1 & biasReg_1[15]) begin // @[BiasActivation.scala 67:85]
        actReg_1 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_1[28] & ~sumReg_1 & ~biasReg_1[15]) begin // @[BiasActivation.scala 70:92]
        actReg_1 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_1 <= _truncWire_1_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_1 <= 16'sh0;
    end
    if ($signed(truncWire_2) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_2[28] & sumReg_2 & biasReg_2[15]) begin // @[BiasActivation.scala 67:85]
        actReg_2 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_2[28] & ~sumReg_2 & ~biasReg_2[15]) begin // @[BiasActivation.scala 70:92]
        actReg_2 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_2 <= _truncWire_2_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_2 <= 16'sh0;
    end
    if ($signed(truncWire_3) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_3[28] & sumReg_3 & biasReg_3[15]) begin // @[BiasActivation.scala 67:85]
        actReg_3 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_3[28] & ~sumReg_3 & ~biasReg_3[15]) begin // @[BiasActivation.scala 70:92]
        actReg_3 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_3 <= _truncWire_3_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_3 <= 16'sh0;
    end
    if ($signed(truncWire_4) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_4[28] & sumReg_4 & biasReg_4[15]) begin // @[BiasActivation.scala 67:85]
        actReg_4 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_4[28] & ~sumReg_4 & ~biasReg_4[15]) begin // @[BiasActivation.scala 70:92]
        actReg_4 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_4 <= _truncWire_4_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_4 <= 16'sh0;
    end
    if ($signed(truncWire_5) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_5[28] & sumReg_5 & biasReg_5[15]) begin // @[BiasActivation.scala 67:85]
        actReg_5 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_5[28] & ~sumReg_5 & ~biasReg_5[15]) begin // @[BiasActivation.scala 70:92]
        actReg_5 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_5 <= _truncWire_5_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_5 <= 16'sh0;
    end
    if ($signed(truncWire_6) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_6[28] & sumReg_6 & biasReg_6[15]) begin // @[BiasActivation.scala 67:85]
        actReg_6 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_6[28] & ~sumReg_6 & ~biasReg_6[15]) begin // @[BiasActivation.scala 70:92]
        actReg_6 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_6 <= _truncWire_6_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_6 <= 16'sh0;
    end
    if ($signed(truncWire_7) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_7[28] & sumReg_7 & biasReg_7[15]) begin // @[BiasActivation.scala 67:85]
        actReg_7 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_7[28] & ~sumReg_7 & ~biasReg_7[15]) begin // @[BiasActivation.scala 70:92]
        actReg_7 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_7 <= _truncWire_7_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_7 <= 16'sh0;
    end
    if ($signed(truncWire_8) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_8[28] & sumReg_8 & biasReg_8[15]) begin // @[BiasActivation.scala 67:85]
        actReg_8 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_8[28] & ~sumReg_8 & ~biasReg_8[15]) begin // @[BiasActivation.scala 70:92]
        actReg_8 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_8 <= _truncWire_8_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_8 <= 16'sh0;
    end
    if ($signed(truncWire_9) >= 16'sh0) begin // @[BiasActivation.scala 80:42]
      if (~plusReg_9[28] & sumReg_9 & biasReg_9[15]) begin // @[BiasActivation.scala 67:85]
        actReg_9 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
      end else if (plusReg_9[28] & ~sumReg_9 & ~biasReg_9[15]) begin // @[BiasActivation.scala 70:92]
        actReg_9 <= 16'sh8000; // @[BiasActivation.scala 72:15]
      end else begin
        actReg_9 <= _truncWire_9_T_1; // @[BiasActivation.scala 74:15]
      end
    end else begin
      actReg_9 <= 16'sh0;
    end
    sumReg_0 <= io_inSum_0[28]; // @[BiasActivation.scala 61:59]
    sumReg_1 <= io_inSum_1[28]; // @[BiasActivation.scala 61:59]
    sumReg_2 <= io_inSum_2[28]; // @[BiasActivation.scala 61:59]
    sumReg_3 <= io_inSum_3[28]; // @[BiasActivation.scala 61:59]
    sumReg_4 <= io_inSum_4[28]; // @[BiasActivation.scala 61:59]
    sumReg_5 <= io_inSum_5[28]; // @[BiasActivation.scala 61:59]
    sumReg_6 <= io_inSum_6[28]; // @[BiasActivation.scala 61:59]
    sumReg_7 <= io_inSum_7[28]; // @[BiasActivation.scala 61:59]
    sumReg_8 <= io_inSum_8[28]; // @[BiasActivation.scala 61:59]
    sumReg_9 <= io_inSum_9[28]; // @[BiasActivation.scala 61:59]
    validReg <= io_inBiasValid; // @[BiasActivation.scala 32:26]
  end
endmodule
module BiasActivation_2(
  input         clock,
  input  [39:0] io_inSum_0,
  input  [39:0] io_inSum_1,
  input  [39:0] io_inSum_2,
  input  [39:0] io_inSum_3,
  input  [39:0] io_inSum_4,
  input  [39:0] io_inSum_5,
  input  [39:0] io_inSum_6,
  input  [39:0] io_inSum_7,
  output [15:0] io_outAct_0,
  output [15:0] io_outAct_1,
  output [15:0] io_outAct_2,
  output [15:0] io_outAct_3,
  output [15:0] io_outAct_4,
  output [15:0] io_outAct_5,
  output [15:0] io_outAct_6,
  output [15:0] io_outAct_7,
  input  [15:0] io_inBias_0,
  input  [15:0] io_inBias_1,
  input  [15:0] io_inBias_2,
  input  [15:0] io_inBias_3,
  input  [15:0] io_inBias_4,
  input  [15:0] io_inBias_5,
  input  [15:0] io_inBias_6,
  input  [15:0] io_inBias_7,
  input         io_inBiasValid
);
  reg [15:0] biasReg_0; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_1; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_2; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_3; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_4; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_5; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_6; // @[BiasActivation.scala 28:22]
  reg [15:0] biasReg_7; // @[BiasActivation.scala 28:22]
  reg [39:0] plusReg_0; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_1; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_2; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_3; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_4; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_5; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_6; // @[BiasActivation.scala 29:22]
  reg [39:0] plusReg_7; // @[BiasActivation.scala 29:22]
  reg [15:0] actReg_0; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_1; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_2; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_3; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_4; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_5; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_6; // @[BiasActivation.scala 30:22]
  reg [15:0] actReg_7; // @[BiasActivation.scala 30:22]
  reg  sumReg_0; // @[BiasActivation.scala 31:22]
  reg  sumReg_1; // @[BiasActivation.scala 31:22]
  reg  sumReg_2; // @[BiasActivation.scala 31:22]
  reg  sumReg_3; // @[BiasActivation.scala 31:22]
  reg  sumReg_4; // @[BiasActivation.scala 31:22]
  reg  sumReg_5; // @[BiasActivation.scala 31:22]
  reg  sumReg_6; // @[BiasActivation.scala 31:22]
  reg  sumReg_7; // @[BiasActivation.scala 31:22]
  reg  validReg; // @[BiasActivation.scala 32:26]
  wire [27:0] _T = {$signed(biasReg_0), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_24 = {{12{_T[27]}},_T}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_4 = {$signed(biasReg_1), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_25 = {{12{_T_4[27]}},_T_4}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_8 = {$signed(biasReg_2), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_26 = {{12{_T_8[27]}},_T_8}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_12 = {$signed(biasReg_3), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_27 = {{12{_T_12[27]}},_T_12}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_16 = {$signed(biasReg_4), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_28 = {{12{_T_16[27]}},_T_16}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_20 = {$signed(biasReg_5), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_29 = {{12{_T_20[27]}},_T_20}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_24 = {$signed(biasReg_6), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_30 = {{12{_T_24[27]}},_T_24}; // @[BiasActivation.scala 56:80]
  wire [27:0] _T_28 = {$signed(biasReg_7), 12'h0}; // @[BiasActivation.scala 56:58]
  wire [39:0] _GEN_31 = {{12{_T_28[27]}},_T_28}; // @[BiasActivation.scala 56:80]
  wire [15:0] _truncWire_0_T_1 = plusReg_0[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_1_T_1 = plusReg_1[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_2_T_1 = plusReg_2[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_3_T_1 = plusReg_3[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_4_T_1 = plusReg_4[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_5_T_1 = plusReg_5[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_6_T_1 = plusReg_6[26:11]; // @[BiasActivation.scala 74:66]
  wire [15:0] _truncWire_7_T_1 = plusReg_7[26:11]; // @[BiasActivation.scala 74:66]
  assign io_outAct_0 = actReg_0; // @[BiasActivation.scala 91:15]
  assign io_outAct_1 = actReg_1; // @[BiasActivation.scala 91:15]
  assign io_outAct_2 = actReg_2; // @[BiasActivation.scala 91:15]
  assign io_outAct_3 = actReg_3; // @[BiasActivation.scala 91:15]
  assign io_outAct_4 = actReg_4; // @[BiasActivation.scala 91:15]
  assign io_outAct_5 = actReg_5; // @[BiasActivation.scala 91:15]
  assign io_outAct_6 = actReg_6; // @[BiasActivation.scala 91:15]
  assign io_outAct_7 = actReg_7; // @[BiasActivation.scala 91:15]
  always @(posedge clock) begin
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_0 <= io_inBias_0; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_1 <= io_inBias_1; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_2 <= io_inBias_2; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_3 <= io_inBias_3; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_4 <= io_inBias_4; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_5 <= io_inBias_5; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_6 <= io_inBias_6; // @[BiasActivation.scala 50:17]
    end
    if (validReg) begin // @[BiasActivation.scala 49:19]
      biasReg_7 <= io_inBias_7; // @[BiasActivation.scala 50:17]
    end
    plusReg_0 <= $signed(_GEN_24) + $signed(io_inSum_0); // @[BiasActivation.scala 56:80]
    plusReg_1 <= $signed(_GEN_25) + $signed(io_inSum_1); // @[BiasActivation.scala 56:80]
    plusReg_2 <= $signed(_GEN_26) + $signed(io_inSum_2); // @[BiasActivation.scala 56:80]
    plusReg_3 <= $signed(_GEN_27) + $signed(io_inSum_3); // @[BiasActivation.scala 56:80]
    plusReg_4 <= $signed(_GEN_28) + $signed(io_inSum_4); // @[BiasActivation.scala 56:80]
    plusReg_5 <= $signed(_GEN_29) + $signed(io_inSum_5); // @[BiasActivation.scala 56:80]
    plusReg_6 <= $signed(_GEN_30) + $signed(io_inSum_6); // @[BiasActivation.scala 56:80]
    plusReg_7 <= $signed(_GEN_31) + $signed(io_inSum_7); // @[BiasActivation.scala 56:80]
    if (~plusReg_0[26] & sumReg_0 & biasReg_0[15]) begin // @[BiasActivation.scala 67:85]
      actReg_0 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_0[26] & ~sumReg_0 & ~biasReg_0[15]) begin // @[BiasActivation.scala 70:92]
      actReg_0 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_0 <= _truncWire_0_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_1[26] & sumReg_1 & biasReg_1[15]) begin // @[BiasActivation.scala 67:85]
      actReg_1 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_1[26] & ~sumReg_1 & ~biasReg_1[15]) begin // @[BiasActivation.scala 70:92]
      actReg_1 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_1 <= _truncWire_1_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_2[26] & sumReg_2 & biasReg_2[15]) begin // @[BiasActivation.scala 67:85]
      actReg_2 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_2[26] & ~sumReg_2 & ~biasReg_2[15]) begin // @[BiasActivation.scala 70:92]
      actReg_2 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_2 <= _truncWire_2_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_3[26] & sumReg_3 & biasReg_3[15]) begin // @[BiasActivation.scala 67:85]
      actReg_3 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_3[26] & ~sumReg_3 & ~biasReg_3[15]) begin // @[BiasActivation.scala 70:92]
      actReg_3 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_3 <= _truncWire_3_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_4[26] & sumReg_4 & biasReg_4[15]) begin // @[BiasActivation.scala 67:85]
      actReg_4 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_4[26] & ~sumReg_4 & ~biasReg_4[15]) begin // @[BiasActivation.scala 70:92]
      actReg_4 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_4 <= _truncWire_4_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_5[26] & sumReg_5 & biasReg_5[15]) begin // @[BiasActivation.scala 67:85]
      actReg_5 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_5[26] & ~sumReg_5 & ~biasReg_5[15]) begin // @[BiasActivation.scala 70:92]
      actReg_5 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_5 <= _truncWire_5_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_6[26] & sumReg_6 & biasReg_6[15]) begin // @[BiasActivation.scala 67:85]
      actReg_6 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_6[26] & ~sumReg_6 & ~biasReg_6[15]) begin // @[BiasActivation.scala 70:92]
      actReg_6 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_6 <= _truncWire_6_T_1; // @[BiasActivation.scala 74:15]
    end
    if (~plusReg_7[26] & sumReg_7 & biasReg_7[15]) begin // @[BiasActivation.scala 67:85]
      actReg_7 <= 16'sh7fff; // @[BiasActivation.scala 69:15]
    end else if (plusReg_7[26] & ~sumReg_7 & ~biasReg_7[15]) begin // @[BiasActivation.scala 70:92]
      actReg_7 <= 16'sh8000; // @[BiasActivation.scala 72:15]
    end else begin
      actReg_7 <= _truncWire_7_T_1; // @[BiasActivation.scala 74:15]
    end
    sumReg_0 <= io_inSum_0[26]; // @[BiasActivation.scala 61:59]
    sumReg_1 <= io_inSum_1[26]; // @[BiasActivation.scala 61:59]
    sumReg_2 <= io_inSum_2[26]; // @[BiasActivation.scala 61:59]
    sumReg_3 <= io_inSum_3[26]; // @[BiasActivation.scala 61:59]
    sumReg_4 <= io_inSum_4[26]; // @[BiasActivation.scala 61:59]
    sumReg_5 <= io_inSum_5[26]; // @[BiasActivation.scala 61:59]
    sumReg_6 <= io_inSum_6[26]; // @[BiasActivation.scala 61:59]
    sumReg_7 <= io_inSum_7[26]; // @[BiasActivation.scala 61:59]
    validReg <= io_inBiasValid; // @[BiasActivation.scala 32:26]
  end
endmodule
module RVTDNN(
  input         clock,
  input  [15:0] io_inAct_0,
  input  [15:0] io_inAct_1,
  input  [15:0] io_inAct_2,
  input  [15:0] io_inAct_3,
  input  [15:0] io_inAct_4,
  input  [15:0] io_inAct_5,
  input  [15:0] io_inAct_6,
  input  [15:0] io_inAct_7,
  output [15:0] io_outAct_0,
  output [15:0] io_outAct_1,
  output [15:0] io_outAct_2,
  output [15:0] io_outAct_3,
  output [15:0] io_outAct_4,
  output [15:0] io_outAct_5,
  output [15:0] io_outAct_6,
  output [15:0] io_outAct_7,
  input  [15:0] io_inWeight_0,
  input  [15:0] io_inWeight_1,
  input  [15:0] io_inWeight_2,
  input  [15:0] io_inWeight_3,
  input  [15:0] io_inWeight_4,
  input  [15:0] io_inWeight_5,
  input  [15:0] io_inWeight_6,
  input  [15:0] io_inWeight_7,
  input  [15:0] io_inWeight_8,
  input  [15:0] io_inWeight_9,
  input  [15:0] io_inBias_0,
  input  [15:0] io_inBias_1,
  input  [15:0] io_inBias_2,
  input  [15:0] io_inBias_3,
  input  [15:0] io_inBias_4,
  input  [15:0] io_inBias_5,
  input  [15:0] io_inBias_6,
  input  [15:0] io_inBias_7,
  input  [15:0] io_inBias_8,
  input  [15:0] io_inBias_9,
  input  [2:0]  io_inWtValid,
  input  [2:0]  io_inBiasValid
);
  wire  SA_0_clock; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_7; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_8; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_9; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_10; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_11; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_12; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_13; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_14; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_15; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_16; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_17; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_18; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inAct_19; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_7; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_8; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_0_io_inWeight_9; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_0; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_1; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_2; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_3; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_4; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_5; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_6; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_7; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_8; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_0_io_outSum_9; // @[RVTDNN.scala 45:48]
  wire  SA_0_io_inwtValid; // @[RVTDNN.scala 45:48]
  wire  SA_1_clock; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_7; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_8; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inAct_9; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_7; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_8; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_1_io_inWeight_9; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_0; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_1; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_2; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_3; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_4; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_5; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_6; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_7; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_8; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_1_io_outSum_9; // @[RVTDNN.scala 45:48]
  wire  SA_1_io_inwtValid; // @[RVTDNN.scala 45:48]
  wire  SA_2_clock; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_7; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_8; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inAct_9; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_0; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_1; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_2; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_3; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_4; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_5; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_6; // @[RVTDNN.scala 45:48]
  wire [15:0] SA_2_io_inWeight_7; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_0; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_1; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_2; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_3; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_4; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_5; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_6; // @[RVTDNN.scala 45:48]
  wire [39:0] SA_2_io_outSum_7; // @[RVTDNN.scala 45:48]
  wire  SA_2_io_inwtValid; // @[RVTDNN.scala 45:48]
  wire  BA_0_clock; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_0; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_1; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_2; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_3; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_4; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_5; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_6; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_7; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_8; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_0_io_inSum_9; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_0; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_1; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_2; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_3; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_4; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_5; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_6; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_7; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_8; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_outAct_9; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_0; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_1; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_2; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_3; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_4; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_5; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_6; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_7; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_8; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_0_io_inBias_9; // @[RVTDNN.scala 52:19]
  wire  BA_0_io_inBiasValid; // @[RVTDNN.scala 52:19]
  wire  BA_1_clock; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_0; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_1; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_2; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_3; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_4; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_5; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_6; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_7; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_8; // @[RVTDNN.scala 52:19]
  wire [39:0] BA_1_io_inSum_9; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_0; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_1; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_2; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_3; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_4; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_5; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_6; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_7; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_8; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_outAct_9; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_0; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_1; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_2; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_3; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_4; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_5; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_6; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_7; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_8; // @[RVTDNN.scala 52:19]
  wire [15:0] BA_1_io_inBias_9; // @[RVTDNN.scala 52:19]
  wire  BA_1_io_inBiasValid; // @[RVTDNN.scala 52:19]
  wire  BA_2_clock; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_0; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_1; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_2; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_3; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_4; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_5; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_6; // @[RVTDNN.scala 48:19]
  wire [39:0] BA_2_io_inSum_7; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_0; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_1; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_2; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_3; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_4; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_5; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_6; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_outAct_7; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_0; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_1; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_2; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_3; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_4; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_5; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_6; // @[RVTDNN.scala 48:19]
  wire [15:0] BA_2_io_inBias_7; // @[RVTDNN.scala 48:19]
  wire  BA_2_io_inBiasValid; // @[RVTDNN.scala 48:19]
  reg [15:0] weightReg_0; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_1; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_2; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_3; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_4; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_5; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_6; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_7; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_8; // @[RVTDNN.scala 28:24]
  reg [15:0] weightReg_9; // @[RVTDNN.scala 28:24]
  reg [15:0] biasReg_0; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_1; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_2; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_3; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_4; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_5; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_6; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_7; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_8; // @[RVTDNN.scala 30:24]
  reg [15:0] biasReg_9; // @[RVTDNN.scala 30:24]
  reg [15:0] inputReg_0_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_1_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_1_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_2_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_2_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_2_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_3_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_3_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_3_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_3_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_4_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_4_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_4_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_4_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_4_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_5_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_6_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_7_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_8_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_9_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_10_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_11_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_12_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_13_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_14_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_15_15; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_15; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_16_16; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_15; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_16; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_17_17; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_15; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_16; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_17; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_18_18; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_0; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_1; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_2; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_3; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_4; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_5; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_6; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_7; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_8; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_9; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_10; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_11; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_12; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_13; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_14; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_15; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_16; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_17; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_18; // @[RVTDNN.scala 36:62]
  reg [15:0] inputReg_19_19; // @[RVTDNN.scala 36:62]
  reg [15:0] outputReg_0_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_1_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_1_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_2_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_2_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_2_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_3_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_3_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_3_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_3_3; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_4_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_4_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_4_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_4_3; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_4_4; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_3; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_4; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_5_5; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_3; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_4; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_5; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_6_6; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_0; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_1; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_2; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_3; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_4; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_5; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_6; // @[RVTDNN.scala 37:62]
  reg [15:0] outputReg_7_7; // @[RVTDNN.scala 37:62]
  wire [159:0] _T_10 = {weightReg_9,weightReg_8,weightReg_7,weightReg_6,weightReg_5,weightReg_4,weightReg_3,weightReg_2,
    weightReg_1,weightReg_0}; // @[RVTDNN.scala 60:59]
  wire [159:0] _T_99 = {biasReg_9,biasReg_8,biasReg_7,biasReg_6,biasReg_5,biasReg_4,biasReg_3,biasReg_2,biasReg_1,
    biasReg_0}; // @[RVTDNN.scala 64:55]
  SystolicArray SA_0 ( // @[RVTDNN.scala 45:48]
    .clock(SA_0_clock),
    .io_inAct_0(SA_0_io_inAct_0),
    .io_inAct_1(SA_0_io_inAct_1),
    .io_inAct_2(SA_0_io_inAct_2),
    .io_inAct_3(SA_0_io_inAct_3),
    .io_inAct_4(SA_0_io_inAct_4),
    .io_inAct_5(SA_0_io_inAct_5),
    .io_inAct_6(SA_0_io_inAct_6),
    .io_inAct_7(SA_0_io_inAct_7),
    .io_inAct_8(SA_0_io_inAct_8),
    .io_inAct_9(SA_0_io_inAct_9),
    .io_inAct_10(SA_0_io_inAct_10),
    .io_inAct_11(SA_0_io_inAct_11),
    .io_inAct_12(SA_0_io_inAct_12),
    .io_inAct_13(SA_0_io_inAct_13),
    .io_inAct_14(SA_0_io_inAct_14),
    .io_inAct_15(SA_0_io_inAct_15),
    .io_inAct_16(SA_0_io_inAct_16),
    .io_inAct_17(SA_0_io_inAct_17),
    .io_inAct_18(SA_0_io_inAct_18),
    .io_inAct_19(SA_0_io_inAct_19),
    .io_inWeight_0(SA_0_io_inWeight_0),
    .io_inWeight_1(SA_0_io_inWeight_1),
    .io_inWeight_2(SA_0_io_inWeight_2),
    .io_inWeight_3(SA_0_io_inWeight_3),
    .io_inWeight_4(SA_0_io_inWeight_4),
    .io_inWeight_5(SA_0_io_inWeight_5),
    .io_inWeight_6(SA_0_io_inWeight_6),
    .io_inWeight_7(SA_0_io_inWeight_7),
    .io_inWeight_8(SA_0_io_inWeight_8),
    .io_inWeight_9(SA_0_io_inWeight_9),
    .io_outSum_0(SA_0_io_outSum_0),
    .io_outSum_1(SA_0_io_outSum_1),
    .io_outSum_2(SA_0_io_outSum_2),
    .io_outSum_3(SA_0_io_outSum_3),
    .io_outSum_4(SA_0_io_outSum_4),
    .io_outSum_5(SA_0_io_outSum_5),
    .io_outSum_6(SA_0_io_outSum_6),
    .io_outSum_7(SA_0_io_outSum_7),
    .io_outSum_8(SA_0_io_outSum_8),
    .io_outSum_9(SA_0_io_outSum_9),
    .io_inwtValid(SA_0_io_inwtValid)
  );
  SystolicArray_1 SA_1 ( // @[RVTDNN.scala 45:48]
    .clock(SA_1_clock),
    .io_inAct_0(SA_1_io_inAct_0),
    .io_inAct_1(SA_1_io_inAct_1),
    .io_inAct_2(SA_1_io_inAct_2),
    .io_inAct_3(SA_1_io_inAct_3),
    .io_inAct_4(SA_1_io_inAct_4),
    .io_inAct_5(SA_1_io_inAct_5),
    .io_inAct_6(SA_1_io_inAct_6),
    .io_inAct_7(SA_1_io_inAct_7),
    .io_inAct_8(SA_1_io_inAct_8),
    .io_inAct_9(SA_1_io_inAct_9),
    .io_inWeight_0(SA_1_io_inWeight_0),
    .io_inWeight_1(SA_1_io_inWeight_1),
    .io_inWeight_2(SA_1_io_inWeight_2),
    .io_inWeight_3(SA_1_io_inWeight_3),
    .io_inWeight_4(SA_1_io_inWeight_4),
    .io_inWeight_5(SA_1_io_inWeight_5),
    .io_inWeight_6(SA_1_io_inWeight_6),
    .io_inWeight_7(SA_1_io_inWeight_7),
    .io_inWeight_8(SA_1_io_inWeight_8),
    .io_inWeight_9(SA_1_io_inWeight_9),
    .io_outSum_0(SA_1_io_outSum_0),
    .io_outSum_1(SA_1_io_outSum_1),
    .io_outSum_2(SA_1_io_outSum_2),
    .io_outSum_3(SA_1_io_outSum_3),
    .io_outSum_4(SA_1_io_outSum_4),
    .io_outSum_5(SA_1_io_outSum_5),
    .io_outSum_6(SA_1_io_outSum_6),
    .io_outSum_7(SA_1_io_outSum_7),
    .io_outSum_8(SA_1_io_outSum_8),
    .io_outSum_9(SA_1_io_outSum_9),
    .io_inwtValid(SA_1_io_inwtValid)
  );
  SystolicArray_2 SA_2 ( // @[RVTDNN.scala 45:48]
    .clock(SA_2_clock),
    .io_inAct_0(SA_2_io_inAct_0),
    .io_inAct_1(SA_2_io_inAct_1),
    .io_inAct_2(SA_2_io_inAct_2),
    .io_inAct_3(SA_2_io_inAct_3),
    .io_inAct_4(SA_2_io_inAct_4),
    .io_inAct_5(SA_2_io_inAct_5),
    .io_inAct_6(SA_2_io_inAct_6),
    .io_inAct_7(SA_2_io_inAct_7),
    .io_inAct_8(SA_2_io_inAct_8),
    .io_inAct_9(SA_2_io_inAct_9),
    .io_inWeight_0(SA_2_io_inWeight_0),
    .io_inWeight_1(SA_2_io_inWeight_1),
    .io_inWeight_2(SA_2_io_inWeight_2),
    .io_inWeight_3(SA_2_io_inWeight_3),
    .io_inWeight_4(SA_2_io_inWeight_4),
    .io_inWeight_5(SA_2_io_inWeight_5),
    .io_inWeight_6(SA_2_io_inWeight_6),
    .io_inWeight_7(SA_2_io_inWeight_7),
    .io_outSum_0(SA_2_io_outSum_0),
    .io_outSum_1(SA_2_io_outSum_1),
    .io_outSum_2(SA_2_io_outSum_2),
    .io_outSum_3(SA_2_io_outSum_3),
    .io_outSum_4(SA_2_io_outSum_4),
    .io_outSum_5(SA_2_io_outSum_5),
    .io_outSum_6(SA_2_io_outSum_6),
    .io_outSum_7(SA_2_io_outSum_7),
    .io_inwtValid(SA_2_io_inwtValid)
  );
  BiasActivation BA_0 ( // @[RVTDNN.scala 52:19]
    .clock(BA_0_clock),
    .io_inSum_0(BA_0_io_inSum_0),
    .io_inSum_1(BA_0_io_inSum_1),
    .io_inSum_2(BA_0_io_inSum_2),
    .io_inSum_3(BA_0_io_inSum_3),
    .io_inSum_4(BA_0_io_inSum_4),
    .io_inSum_5(BA_0_io_inSum_5),
    .io_inSum_6(BA_0_io_inSum_6),
    .io_inSum_7(BA_0_io_inSum_7),
    .io_inSum_8(BA_0_io_inSum_8),
    .io_inSum_9(BA_0_io_inSum_9),
    .io_outAct_0(BA_0_io_outAct_0),
    .io_outAct_1(BA_0_io_outAct_1),
    .io_outAct_2(BA_0_io_outAct_2),
    .io_outAct_3(BA_0_io_outAct_3),
    .io_outAct_4(BA_0_io_outAct_4),
    .io_outAct_5(BA_0_io_outAct_5),
    .io_outAct_6(BA_0_io_outAct_6),
    .io_outAct_7(BA_0_io_outAct_7),
    .io_outAct_8(BA_0_io_outAct_8),
    .io_outAct_9(BA_0_io_outAct_9),
    .io_inBias_0(BA_0_io_inBias_0),
    .io_inBias_1(BA_0_io_inBias_1),
    .io_inBias_2(BA_0_io_inBias_2),
    .io_inBias_3(BA_0_io_inBias_3),
    .io_inBias_4(BA_0_io_inBias_4),
    .io_inBias_5(BA_0_io_inBias_5),
    .io_inBias_6(BA_0_io_inBias_6),
    .io_inBias_7(BA_0_io_inBias_7),
    .io_inBias_8(BA_0_io_inBias_8),
    .io_inBias_9(BA_0_io_inBias_9),
    .io_inBiasValid(BA_0_io_inBiasValid)
  );
  BiasActivation_1 BA_1 ( // @[RVTDNN.scala 52:19]
    .clock(BA_1_clock),
    .io_inSum_0(BA_1_io_inSum_0),
    .io_inSum_1(BA_1_io_inSum_1),
    .io_inSum_2(BA_1_io_inSum_2),
    .io_inSum_3(BA_1_io_inSum_3),
    .io_inSum_4(BA_1_io_inSum_4),
    .io_inSum_5(BA_1_io_inSum_5),
    .io_inSum_6(BA_1_io_inSum_6),
    .io_inSum_7(BA_1_io_inSum_7),
    .io_inSum_8(BA_1_io_inSum_8),
    .io_inSum_9(BA_1_io_inSum_9),
    .io_outAct_0(BA_1_io_outAct_0),
    .io_outAct_1(BA_1_io_outAct_1),
    .io_outAct_2(BA_1_io_outAct_2),
    .io_outAct_3(BA_1_io_outAct_3),
    .io_outAct_4(BA_1_io_outAct_4),
    .io_outAct_5(BA_1_io_outAct_5),
    .io_outAct_6(BA_1_io_outAct_6),
    .io_outAct_7(BA_1_io_outAct_7),
    .io_outAct_8(BA_1_io_outAct_8),
    .io_outAct_9(BA_1_io_outAct_9),
    .io_inBias_0(BA_1_io_inBias_0),
    .io_inBias_1(BA_1_io_inBias_1),
    .io_inBias_2(BA_1_io_inBias_2),
    .io_inBias_3(BA_1_io_inBias_3),
    .io_inBias_4(BA_1_io_inBias_4),
    .io_inBias_5(BA_1_io_inBias_5),
    .io_inBias_6(BA_1_io_inBias_6),
    .io_inBias_7(BA_1_io_inBias_7),
    .io_inBias_8(BA_1_io_inBias_8),
    .io_inBias_9(BA_1_io_inBias_9),
    .io_inBiasValid(BA_1_io_inBiasValid)
  );
  BiasActivation_2 BA_2 ( // @[RVTDNN.scala 48:19]
    .clock(BA_2_clock),
    .io_inSum_0(BA_2_io_inSum_0),
    .io_inSum_1(BA_2_io_inSum_1),
    .io_inSum_2(BA_2_io_inSum_2),
    .io_inSum_3(BA_2_io_inSum_3),
    .io_inSum_4(BA_2_io_inSum_4),
    .io_inSum_5(BA_2_io_inSum_5),
    .io_inSum_6(BA_2_io_inSum_6),
    .io_inSum_7(BA_2_io_inSum_7),
    .io_outAct_0(BA_2_io_outAct_0),
    .io_outAct_1(BA_2_io_outAct_1),
    .io_outAct_2(BA_2_io_outAct_2),
    .io_outAct_3(BA_2_io_outAct_3),
    .io_outAct_4(BA_2_io_outAct_4),
    .io_outAct_5(BA_2_io_outAct_5),
    .io_outAct_6(BA_2_io_outAct_6),
    .io_outAct_7(BA_2_io_outAct_7),
    .io_inBias_0(BA_2_io_inBias_0),
    .io_inBias_1(BA_2_io_inBias_1),
    .io_inBias_2(BA_2_io_inBias_2),
    .io_inBias_3(BA_2_io_inBias_3),
    .io_inBias_4(BA_2_io_inBias_4),
    .io_inBias_5(BA_2_io_inBias_5),
    .io_inBias_6(BA_2_io_inBias_6),
    .io_inBias_7(BA_2_io_inBias_7),
    .io_inBiasValid(BA_2_io_inBiasValid)
  );
  assign io_outAct_0 = outputReg_0_0; // @[RVTDNN.scala 75:15]
  assign io_outAct_1 = outputReg_1_1; // @[RVTDNN.scala 75:15]
  assign io_outAct_2 = outputReg_2_2; // @[RVTDNN.scala 75:15]
  assign io_outAct_3 = outputReg_3_3; // @[RVTDNN.scala 75:15]
  assign io_outAct_4 = outputReg_4_4; // @[RVTDNN.scala 75:15]
  assign io_outAct_5 = outputReg_5_5; // @[RVTDNN.scala 75:15]
  assign io_outAct_6 = outputReg_6_6; // @[RVTDNN.scala 75:15]
  assign io_outAct_7 = outputReg_7_7; // @[RVTDNN.scala 75:15]
  assign SA_0_clock = clock;
  assign SA_0_io_inAct_0 = inputReg_0_0; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_1 = inputReg_1_1; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_2 = inputReg_2_2; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_3 = inputReg_3_3; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_4 = inputReg_4_4; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_5 = inputReg_5_5; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_6 = inputReg_6_6; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_7 = inputReg_7_7; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_8 = inputReg_8_8; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_9 = inputReg_9_9; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_10 = inputReg_10_10; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_11 = inputReg_11_11; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_12 = inputReg_12_12; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_13 = inputReg_13_13; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_14 = inputReg_14_14; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_15 = inputReg_15_15; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_16 = inputReg_16_16; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_17 = inputReg_17_17; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_18 = inputReg_18_18; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inAct_19 = inputReg_19_19; // @[RVTDNN.scala 79:35]
  assign SA_0_io_inWeight_0 = _T_10[15:0]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_1 = _T_10[31:16]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_2 = _T_10[47:32]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_3 = _T_10[63:48]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_4 = _T_10[79:64]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_5 = _T_10[95:80]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_6 = _T_10[111:96]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_7 = _T_10[127:112]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_8 = _T_10[143:128]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inWeight_9 = _T_10[159:144]; // @[RVTDNN.scala 60:59]
  assign SA_0_io_inwtValid = io_inWtValid[0]; // @[RVTDNN.scala 62:26]
  assign SA_1_clock = clock;
  assign SA_1_io_inAct_0 = BA_0_io_outAct_0; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_1 = BA_0_io_outAct_1; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_2 = BA_0_io_outAct_2; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_3 = BA_0_io_outAct_3; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_4 = BA_0_io_outAct_4; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_5 = BA_0_io_outAct_5; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_6 = BA_0_io_outAct_6; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_7 = BA_0_io_outAct_7; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_8 = BA_0_io_outAct_8; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inAct_9 = BA_0_io_outAct_9; // @[RVTDNN.scala 80:35]
  assign SA_1_io_inWeight_0 = _T_10[15:0]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_1 = _T_10[31:16]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_2 = _T_10[47:32]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_3 = _T_10[63:48]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_4 = _T_10[79:64]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_5 = _T_10[95:80]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_6 = _T_10[111:96]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_7 = _T_10[127:112]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_8 = _T_10[143:128]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inWeight_9 = _T_10[159:144]; // @[RVTDNN.scala 60:59]
  assign SA_1_io_inwtValid = io_inWtValid[1]; // @[RVTDNN.scala 62:26]
  assign SA_2_clock = clock;
  assign SA_2_io_inAct_0 = BA_1_io_outAct_0; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_1 = BA_1_io_outAct_1; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_2 = BA_1_io_outAct_2; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_3 = BA_1_io_outAct_3; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_4 = BA_1_io_outAct_4; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_5 = BA_1_io_outAct_5; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_6 = BA_1_io_outAct_6; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_7 = BA_1_io_outAct_7; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_8 = BA_1_io_outAct_8; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inAct_9 = BA_1_io_outAct_9; // @[RVTDNN.scala 80:35]
  assign SA_2_io_inWeight_0 = _T_10[15:0]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_1 = _T_10[31:16]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_2 = _T_10[47:32]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_3 = _T_10[63:48]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_4 = _T_10[79:64]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_5 = _T_10[95:80]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_6 = _T_10[111:96]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inWeight_7 = _T_10[127:112]; // @[RVTDNN.scala 60:59]
  assign SA_2_io_inwtValid = io_inWtValid[2]; // @[RVTDNN.scala 62:26]
  assign BA_0_clock = clock;
  assign BA_0_io_inSum_0 = SA_0_io_outSum_0; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_1 = SA_0_io_outSum_1; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_2 = SA_0_io_outSum_2; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_3 = SA_0_io_outSum_3; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_4 = SA_0_io_outSum_4; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_5 = SA_0_io_outSum_5; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_6 = SA_0_io_outSum_6; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_7 = SA_0_io_outSum_7; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_8 = SA_0_io_outSum_8; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inSum_9 = SA_0_io_outSum_9; // @[RVTDNN.scala 81:24]
  assign BA_0_io_inBias_0 = _T_99[15:0]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_1 = _T_99[31:16]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_2 = _T_99[47:32]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_3 = _T_99[63:48]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_4 = _T_99[79:64]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_5 = _T_99[95:80]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_6 = _T_99[111:96]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_7 = _T_99[127:112]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_8 = _T_99[143:128]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBias_9 = _T_99[159:144]; // @[RVTDNN.scala 64:55]
  assign BA_0_io_inBiasValid = io_inBiasValid[0]; // @[RVTDNN.scala 66:28]
  assign BA_1_clock = clock;
  assign BA_1_io_inSum_0 = SA_1_io_outSum_0; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_1 = SA_1_io_outSum_1; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_2 = SA_1_io_outSum_2; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_3 = SA_1_io_outSum_3; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_4 = SA_1_io_outSum_4; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_5 = SA_1_io_outSum_5; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_6 = SA_1_io_outSum_6; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_7 = SA_1_io_outSum_7; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_8 = SA_1_io_outSum_8; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inSum_9 = SA_1_io_outSum_9; // @[RVTDNN.scala 81:24]
  assign BA_1_io_inBias_0 = _T_99[15:0]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_1 = _T_99[31:16]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_2 = _T_99[47:32]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_3 = _T_99[63:48]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_4 = _T_99[79:64]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_5 = _T_99[95:80]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_6 = _T_99[111:96]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_7 = _T_99[127:112]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_8 = _T_99[143:128]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBias_9 = _T_99[159:144]; // @[RVTDNN.scala 64:55]
  assign BA_1_io_inBiasValid = io_inBiasValid[1]; // @[RVTDNN.scala 66:28]
  assign BA_2_clock = clock;
  assign BA_2_io_inSum_0 = SA_2_io_outSum_0; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_1 = SA_2_io_outSum_1; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_2 = SA_2_io_outSum_2; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_3 = SA_2_io_outSum_3; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_4 = SA_2_io_outSum_4; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_5 = SA_2_io_outSum_5; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_6 = SA_2_io_outSum_6; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inSum_7 = SA_2_io_outSum_7; // @[RVTDNN.scala 81:24]
  assign BA_2_io_inBias_0 = _T_99[15:0]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_1 = _T_99[31:16]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_2 = _T_99[47:32]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_3 = _T_99[63:48]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_4 = _T_99[79:64]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_5 = _T_99[95:80]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_6 = _T_99[111:96]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBias_7 = _T_99[127:112]; // @[RVTDNN.scala 64:55]
  assign BA_2_io_inBiasValid = io_inBiasValid[2]; // @[RVTDNN.scala 66:28]
  always @(posedge clock) begin
    weightReg_0 <= io_inWeight_0; // @[RVTDNN.scala 29:17]
    weightReg_1 <= io_inWeight_1; // @[RVTDNN.scala 29:17]
    weightReg_2 <= io_inWeight_2; // @[RVTDNN.scala 29:17]
    weightReg_3 <= io_inWeight_3; // @[RVTDNN.scala 29:17]
    weightReg_4 <= io_inWeight_4; // @[RVTDNN.scala 29:17]
    weightReg_5 <= io_inWeight_5; // @[RVTDNN.scala 29:17]
    weightReg_6 <= io_inWeight_6; // @[RVTDNN.scala 29:17]
    weightReg_7 <= io_inWeight_7; // @[RVTDNN.scala 29:17]
    weightReg_8 <= io_inWeight_8; // @[RVTDNN.scala 29:17]
    weightReg_9 <= io_inWeight_9; // @[RVTDNN.scala 29:17]
    biasReg_0 <= io_inBias_0; // @[RVTDNN.scala 31:17]
    biasReg_1 <= io_inBias_1; // @[RVTDNN.scala 31:17]
    biasReg_2 <= io_inBias_2; // @[RVTDNN.scala 31:17]
    biasReg_3 <= io_inBias_3; // @[RVTDNN.scala 31:17]
    biasReg_4 <= io_inBias_4; // @[RVTDNN.scala 31:17]
    biasReg_5 <= io_inBias_5; // @[RVTDNN.scala 31:17]
    biasReg_6 <= io_inBias_6; // @[RVTDNN.scala 31:17]
    biasReg_7 <= io_inBias_7; // @[RVTDNN.scala 31:17]
    biasReg_8 <= io_inBias_8; // @[RVTDNN.scala 31:17]
    biasReg_9 <= io_inBias_9; // @[RVTDNN.scala 31:17]
    inputReg_0_0 <= io_inAct_0; // @[RVTDNN.scala 40:25 41:62]
    inputReg_1_0 <= io_inAct_1; // @[RVTDNN.scala 40:25 41:62]
    inputReg_1_1 <= inputReg_1_0; // @[RVTDNN.scala 70:62]
    inputReg_2_0 <= io_inAct_2; // @[RVTDNN.scala 40:25 41:62]
    inputReg_2_1 <= inputReg_2_0; // @[RVTDNN.scala 70:62]
    inputReg_2_2 <= inputReg_2_1; // @[RVTDNN.scala 70:62]
    inputReg_3_0 <= io_inAct_3; // @[RVTDNN.scala 40:25 41:62]
    inputReg_3_1 <= inputReg_3_0; // @[RVTDNN.scala 70:62]
    inputReg_3_2 <= inputReg_3_1; // @[RVTDNN.scala 70:62]
    inputReg_3_3 <= inputReg_3_2; // @[RVTDNN.scala 70:62]
    inputReg_4_0 <= io_inAct_4; // @[RVTDNN.scala 40:25 41:62]
    inputReg_4_1 <= inputReg_4_0; // @[RVTDNN.scala 70:62]
    inputReg_4_2 <= inputReg_4_1; // @[RVTDNN.scala 70:62]
    inputReg_4_3 <= inputReg_4_2; // @[RVTDNN.scala 70:62]
    inputReg_4_4 <= inputReg_4_3; // @[RVTDNN.scala 70:62]
    inputReg_5_0 <= io_inAct_5; // @[RVTDNN.scala 40:25 41:62]
    inputReg_5_1 <= inputReg_5_0; // @[RVTDNN.scala 70:62]
    inputReg_5_2 <= inputReg_5_1; // @[RVTDNN.scala 70:62]
    inputReg_5_3 <= inputReg_5_2; // @[RVTDNN.scala 70:62]
    inputReg_5_4 <= inputReg_5_3; // @[RVTDNN.scala 70:62]
    inputReg_5_5 <= inputReg_5_4; // @[RVTDNN.scala 70:62]
    inputReg_6_0 <= io_inAct_6; // @[RVTDNN.scala 40:25 41:62]
    inputReg_6_1 <= inputReg_6_0; // @[RVTDNN.scala 70:62]
    inputReg_6_2 <= inputReg_6_1; // @[RVTDNN.scala 70:62]
    inputReg_6_3 <= inputReg_6_2; // @[RVTDNN.scala 70:62]
    inputReg_6_4 <= inputReg_6_3; // @[RVTDNN.scala 70:62]
    inputReg_6_5 <= inputReg_6_4; // @[RVTDNN.scala 70:62]
    inputReg_6_6 <= inputReg_6_5; // @[RVTDNN.scala 70:62]
    inputReg_7_0 <= io_inAct_7; // @[RVTDNN.scala 40:25 41:62]
    inputReg_7_1 <= inputReg_7_0; // @[RVTDNN.scala 70:62]
    inputReg_7_2 <= inputReg_7_1; // @[RVTDNN.scala 70:62]
    inputReg_7_3 <= inputReg_7_2; // @[RVTDNN.scala 70:62]
    inputReg_7_4 <= inputReg_7_3; // @[RVTDNN.scala 70:62]
    inputReg_7_5 <= inputReg_7_4; // @[RVTDNN.scala 70:62]
    inputReg_7_6 <= inputReg_7_5; // @[RVTDNN.scala 70:62]
    inputReg_7_7 <= inputReg_7_6; // @[RVTDNN.scala 70:62]
    inputReg_8_0 <= inputReg_0_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_8_1 <= inputReg_8_0; // @[RVTDNN.scala 70:62]
    inputReg_8_2 <= inputReg_8_1; // @[RVTDNN.scala 70:62]
    inputReg_8_3 <= inputReg_8_2; // @[RVTDNN.scala 70:62]
    inputReg_8_4 <= inputReg_8_3; // @[RVTDNN.scala 70:62]
    inputReg_8_5 <= inputReg_8_4; // @[RVTDNN.scala 70:62]
    inputReg_8_6 <= inputReg_8_5; // @[RVTDNN.scala 70:62]
    inputReg_8_7 <= inputReg_8_6; // @[RVTDNN.scala 70:62]
    inputReg_8_8 <= inputReg_8_7; // @[RVTDNN.scala 70:62]
    inputReg_9_0 <= inputReg_1_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_9_1 <= inputReg_9_0; // @[RVTDNN.scala 70:62]
    inputReg_9_2 <= inputReg_9_1; // @[RVTDNN.scala 70:62]
    inputReg_9_3 <= inputReg_9_2; // @[RVTDNN.scala 70:62]
    inputReg_9_4 <= inputReg_9_3; // @[RVTDNN.scala 70:62]
    inputReg_9_5 <= inputReg_9_4; // @[RVTDNN.scala 70:62]
    inputReg_9_6 <= inputReg_9_5; // @[RVTDNN.scala 70:62]
    inputReg_9_7 <= inputReg_9_6; // @[RVTDNN.scala 70:62]
    inputReg_9_8 <= inputReg_9_7; // @[RVTDNN.scala 70:62]
    inputReg_9_9 <= inputReg_9_8; // @[RVTDNN.scala 70:62]
    inputReg_10_0 <= inputReg_2_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_10_1 <= inputReg_10_0; // @[RVTDNN.scala 70:62]
    inputReg_10_2 <= inputReg_10_1; // @[RVTDNN.scala 70:62]
    inputReg_10_3 <= inputReg_10_2; // @[RVTDNN.scala 70:62]
    inputReg_10_4 <= inputReg_10_3; // @[RVTDNN.scala 70:62]
    inputReg_10_5 <= inputReg_10_4; // @[RVTDNN.scala 70:62]
    inputReg_10_6 <= inputReg_10_5; // @[RVTDNN.scala 70:62]
    inputReg_10_7 <= inputReg_10_6; // @[RVTDNN.scala 70:62]
    inputReg_10_8 <= inputReg_10_7; // @[RVTDNN.scala 70:62]
    inputReg_10_9 <= inputReg_10_8; // @[RVTDNN.scala 70:62]
    inputReg_10_10 <= inputReg_10_9; // @[RVTDNN.scala 70:62]
    inputReg_11_0 <= inputReg_3_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_11_1 <= inputReg_11_0; // @[RVTDNN.scala 70:62]
    inputReg_11_2 <= inputReg_11_1; // @[RVTDNN.scala 70:62]
    inputReg_11_3 <= inputReg_11_2; // @[RVTDNN.scala 70:62]
    inputReg_11_4 <= inputReg_11_3; // @[RVTDNN.scala 70:62]
    inputReg_11_5 <= inputReg_11_4; // @[RVTDNN.scala 70:62]
    inputReg_11_6 <= inputReg_11_5; // @[RVTDNN.scala 70:62]
    inputReg_11_7 <= inputReg_11_6; // @[RVTDNN.scala 70:62]
    inputReg_11_8 <= inputReg_11_7; // @[RVTDNN.scala 70:62]
    inputReg_11_9 <= inputReg_11_8; // @[RVTDNN.scala 70:62]
    inputReg_11_10 <= inputReg_11_9; // @[RVTDNN.scala 70:62]
    inputReg_11_11 <= inputReg_11_10; // @[RVTDNN.scala 70:62]
    inputReg_12_0 <= inputReg_4_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_12_1 <= inputReg_12_0; // @[RVTDNN.scala 70:62]
    inputReg_12_2 <= inputReg_12_1; // @[RVTDNN.scala 70:62]
    inputReg_12_3 <= inputReg_12_2; // @[RVTDNN.scala 70:62]
    inputReg_12_4 <= inputReg_12_3; // @[RVTDNN.scala 70:62]
    inputReg_12_5 <= inputReg_12_4; // @[RVTDNN.scala 70:62]
    inputReg_12_6 <= inputReg_12_5; // @[RVTDNN.scala 70:62]
    inputReg_12_7 <= inputReg_12_6; // @[RVTDNN.scala 70:62]
    inputReg_12_8 <= inputReg_12_7; // @[RVTDNN.scala 70:62]
    inputReg_12_9 <= inputReg_12_8; // @[RVTDNN.scala 70:62]
    inputReg_12_10 <= inputReg_12_9; // @[RVTDNN.scala 70:62]
    inputReg_12_11 <= inputReg_12_10; // @[RVTDNN.scala 70:62]
    inputReg_12_12 <= inputReg_12_11; // @[RVTDNN.scala 70:62]
    inputReg_13_0 <= inputReg_5_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_13_1 <= inputReg_13_0; // @[RVTDNN.scala 70:62]
    inputReg_13_2 <= inputReg_13_1; // @[RVTDNN.scala 70:62]
    inputReg_13_3 <= inputReg_13_2; // @[RVTDNN.scala 70:62]
    inputReg_13_4 <= inputReg_13_3; // @[RVTDNN.scala 70:62]
    inputReg_13_5 <= inputReg_13_4; // @[RVTDNN.scala 70:62]
    inputReg_13_6 <= inputReg_13_5; // @[RVTDNN.scala 70:62]
    inputReg_13_7 <= inputReg_13_6; // @[RVTDNN.scala 70:62]
    inputReg_13_8 <= inputReg_13_7; // @[RVTDNN.scala 70:62]
    inputReg_13_9 <= inputReg_13_8; // @[RVTDNN.scala 70:62]
    inputReg_13_10 <= inputReg_13_9; // @[RVTDNN.scala 70:62]
    inputReg_13_11 <= inputReg_13_10; // @[RVTDNN.scala 70:62]
    inputReg_13_12 <= inputReg_13_11; // @[RVTDNN.scala 70:62]
    inputReg_13_13 <= inputReg_13_12; // @[RVTDNN.scala 70:62]
    inputReg_14_0 <= inputReg_6_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_14_1 <= inputReg_14_0; // @[RVTDNN.scala 70:62]
    inputReg_14_2 <= inputReg_14_1; // @[RVTDNN.scala 70:62]
    inputReg_14_3 <= inputReg_14_2; // @[RVTDNN.scala 70:62]
    inputReg_14_4 <= inputReg_14_3; // @[RVTDNN.scala 70:62]
    inputReg_14_5 <= inputReg_14_4; // @[RVTDNN.scala 70:62]
    inputReg_14_6 <= inputReg_14_5; // @[RVTDNN.scala 70:62]
    inputReg_14_7 <= inputReg_14_6; // @[RVTDNN.scala 70:62]
    inputReg_14_8 <= inputReg_14_7; // @[RVTDNN.scala 70:62]
    inputReg_14_9 <= inputReg_14_8; // @[RVTDNN.scala 70:62]
    inputReg_14_10 <= inputReg_14_9; // @[RVTDNN.scala 70:62]
    inputReg_14_11 <= inputReg_14_10; // @[RVTDNN.scala 70:62]
    inputReg_14_12 <= inputReg_14_11; // @[RVTDNN.scala 70:62]
    inputReg_14_13 <= inputReg_14_12; // @[RVTDNN.scala 70:62]
    inputReg_14_14 <= inputReg_14_13; // @[RVTDNN.scala 70:62]
    inputReg_15_0 <= inputReg_7_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_15_1 <= inputReg_15_0; // @[RVTDNN.scala 70:62]
    inputReg_15_2 <= inputReg_15_1; // @[RVTDNN.scala 70:62]
    inputReg_15_3 <= inputReg_15_2; // @[RVTDNN.scala 70:62]
    inputReg_15_4 <= inputReg_15_3; // @[RVTDNN.scala 70:62]
    inputReg_15_5 <= inputReg_15_4; // @[RVTDNN.scala 70:62]
    inputReg_15_6 <= inputReg_15_5; // @[RVTDNN.scala 70:62]
    inputReg_15_7 <= inputReg_15_6; // @[RVTDNN.scala 70:62]
    inputReg_15_8 <= inputReg_15_7; // @[RVTDNN.scala 70:62]
    inputReg_15_9 <= inputReg_15_8; // @[RVTDNN.scala 70:62]
    inputReg_15_10 <= inputReg_15_9; // @[RVTDNN.scala 70:62]
    inputReg_15_11 <= inputReg_15_10; // @[RVTDNN.scala 70:62]
    inputReg_15_12 <= inputReg_15_11; // @[RVTDNN.scala 70:62]
    inputReg_15_13 <= inputReg_15_12; // @[RVTDNN.scala 70:62]
    inputReg_15_14 <= inputReg_15_13; // @[RVTDNN.scala 70:62]
    inputReg_15_15 <= inputReg_15_14; // @[RVTDNN.scala 70:62]
    inputReg_16_0 <= inputReg_8_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_16_1 <= inputReg_16_0; // @[RVTDNN.scala 70:62]
    inputReg_16_2 <= inputReg_16_1; // @[RVTDNN.scala 70:62]
    inputReg_16_3 <= inputReg_16_2; // @[RVTDNN.scala 70:62]
    inputReg_16_4 <= inputReg_16_3; // @[RVTDNN.scala 70:62]
    inputReg_16_5 <= inputReg_16_4; // @[RVTDNN.scala 70:62]
    inputReg_16_6 <= inputReg_16_5; // @[RVTDNN.scala 70:62]
    inputReg_16_7 <= inputReg_16_6; // @[RVTDNN.scala 70:62]
    inputReg_16_8 <= inputReg_16_7; // @[RVTDNN.scala 70:62]
    inputReg_16_9 <= inputReg_16_8; // @[RVTDNN.scala 70:62]
    inputReg_16_10 <= inputReg_16_9; // @[RVTDNN.scala 70:62]
    inputReg_16_11 <= inputReg_16_10; // @[RVTDNN.scala 70:62]
    inputReg_16_12 <= inputReg_16_11; // @[RVTDNN.scala 70:62]
    inputReg_16_13 <= inputReg_16_12; // @[RVTDNN.scala 70:62]
    inputReg_16_14 <= inputReg_16_13; // @[RVTDNN.scala 70:62]
    inputReg_16_15 <= inputReg_16_14; // @[RVTDNN.scala 70:62]
    inputReg_16_16 <= inputReg_16_15; // @[RVTDNN.scala 70:62]
    inputReg_17_0 <= inputReg_9_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_17_1 <= inputReg_17_0; // @[RVTDNN.scala 70:62]
    inputReg_17_2 <= inputReg_17_1; // @[RVTDNN.scala 70:62]
    inputReg_17_3 <= inputReg_17_2; // @[RVTDNN.scala 70:62]
    inputReg_17_4 <= inputReg_17_3; // @[RVTDNN.scala 70:62]
    inputReg_17_5 <= inputReg_17_4; // @[RVTDNN.scala 70:62]
    inputReg_17_6 <= inputReg_17_5; // @[RVTDNN.scala 70:62]
    inputReg_17_7 <= inputReg_17_6; // @[RVTDNN.scala 70:62]
    inputReg_17_8 <= inputReg_17_7; // @[RVTDNN.scala 70:62]
    inputReg_17_9 <= inputReg_17_8; // @[RVTDNN.scala 70:62]
    inputReg_17_10 <= inputReg_17_9; // @[RVTDNN.scala 70:62]
    inputReg_17_11 <= inputReg_17_10; // @[RVTDNN.scala 70:62]
    inputReg_17_12 <= inputReg_17_11; // @[RVTDNN.scala 70:62]
    inputReg_17_13 <= inputReg_17_12; // @[RVTDNN.scala 70:62]
    inputReg_17_14 <= inputReg_17_13; // @[RVTDNN.scala 70:62]
    inputReg_17_15 <= inputReg_17_14; // @[RVTDNN.scala 70:62]
    inputReg_17_16 <= inputReg_17_15; // @[RVTDNN.scala 70:62]
    inputReg_17_17 <= inputReg_17_16; // @[RVTDNN.scala 70:62]
    inputReg_18_0 <= inputReg_10_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_18_1 <= inputReg_18_0; // @[RVTDNN.scala 70:62]
    inputReg_18_2 <= inputReg_18_1; // @[RVTDNN.scala 70:62]
    inputReg_18_3 <= inputReg_18_2; // @[RVTDNN.scala 70:62]
    inputReg_18_4 <= inputReg_18_3; // @[RVTDNN.scala 70:62]
    inputReg_18_5 <= inputReg_18_4; // @[RVTDNN.scala 70:62]
    inputReg_18_6 <= inputReg_18_5; // @[RVTDNN.scala 70:62]
    inputReg_18_7 <= inputReg_18_6; // @[RVTDNN.scala 70:62]
    inputReg_18_8 <= inputReg_18_7; // @[RVTDNN.scala 70:62]
    inputReg_18_9 <= inputReg_18_8; // @[RVTDNN.scala 70:62]
    inputReg_18_10 <= inputReg_18_9; // @[RVTDNN.scala 70:62]
    inputReg_18_11 <= inputReg_18_10; // @[RVTDNN.scala 70:62]
    inputReg_18_12 <= inputReg_18_11; // @[RVTDNN.scala 70:62]
    inputReg_18_13 <= inputReg_18_12; // @[RVTDNN.scala 70:62]
    inputReg_18_14 <= inputReg_18_13; // @[RVTDNN.scala 70:62]
    inputReg_18_15 <= inputReg_18_14; // @[RVTDNN.scala 70:62]
    inputReg_18_16 <= inputReg_18_15; // @[RVTDNN.scala 70:62]
    inputReg_18_17 <= inputReg_18_16; // @[RVTDNN.scala 70:62]
    inputReg_18_18 <= inputReg_18_17; // @[RVTDNN.scala 70:62]
    inputReg_19_0 <= inputReg_11_0; // @[RVTDNN.scala 40:25 42:62]
    inputReg_19_1 <= inputReg_19_0; // @[RVTDNN.scala 70:62]
    inputReg_19_2 <= inputReg_19_1; // @[RVTDNN.scala 70:62]
    inputReg_19_3 <= inputReg_19_2; // @[RVTDNN.scala 70:62]
    inputReg_19_4 <= inputReg_19_3; // @[RVTDNN.scala 70:62]
    inputReg_19_5 <= inputReg_19_4; // @[RVTDNN.scala 70:62]
    inputReg_19_6 <= inputReg_19_5; // @[RVTDNN.scala 70:62]
    inputReg_19_7 <= inputReg_19_6; // @[RVTDNN.scala 70:62]
    inputReg_19_8 <= inputReg_19_7; // @[RVTDNN.scala 70:62]
    inputReg_19_9 <= inputReg_19_8; // @[RVTDNN.scala 70:62]
    inputReg_19_10 <= inputReg_19_9; // @[RVTDNN.scala 70:62]
    inputReg_19_11 <= inputReg_19_10; // @[RVTDNN.scala 70:62]
    inputReg_19_12 <= inputReg_19_11; // @[RVTDNN.scala 70:62]
    inputReg_19_13 <= inputReg_19_12; // @[RVTDNN.scala 70:62]
    inputReg_19_14 <= inputReg_19_13; // @[RVTDNN.scala 70:62]
    inputReg_19_15 <= inputReg_19_14; // @[RVTDNN.scala 70:62]
    inputReg_19_16 <= inputReg_19_15; // @[RVTDNN.scala 70:62]
    inputReg_19_17 <= inputReg_19_16; // @[RVTDNN.scala 70:62]
    inputReg_19_18 <= inputReg_19_17; // @[RVTDNN.scala 70:62]
    inputReg_19_19 <= inputReg_19_18; // @[RVTDNN.scala 70:62]
    outputReg_0_0 <= BA_2_io_outAct_7; // @[RVTDNN.scala 73:63]
    outputReg_1_0 <= BA_2_io_outAct_6; // @[RVTDNN.scala 73:63]
    outputReg_1_1 <= outputReg_1_0; // @[RVTDNN.scala 72:63]
    outputReg_2_0 <= BA_2_io_outAct_5; // @[RVTDNN.scala 73:63]
    outputReg_2_1 <= outputReg_2_0; // @[RVTDNN.scala 72:63]
    outputReg_2_2 <= outputReg_2_1; // @[RVTDNN.scala 72:63]
    outputReg_3_0 <= BA_2_io_outAct_4; // @[RVTDNN.scala 73:63]
    outputReg_3_1 <= outputReg_3_0; // @[RVTDNN.scala 72:63]
    outputReg_3_2 <= outputReg_3_1; // @[RVTDNN.scala 72:63]
    outputReg_3_3 <= outputReg_3_2; // @[RVTDNN.scala 72:63]
    outputReg_4_0 <= BA_2_io_outAct_3; // @[RVTDNN.scala 73:63]
    outputReg_4_1 <= outputReg_4_0; // @[RVTDNN.scala 72:63]
    outputReg_4_2 <= outputReg_4_1; // @[RVTDNN.scala 72:63]
    outputReg_4_3 <= outputReg_4_2; // @[RVTDNN.scala 72:63]
    outputReg_4_4 <= outputReg_4_3; // @[RVTDNN.scala 72:63]
    outputReg_5_0 <= BA_2_io_outAct_2; // @[RVTDNN.scala 73:63]
    outputReg_5_1 <= outputReg_5_0; // @[RVTDNN.scala 72:63]
    outputReg_5_2 <= outputReg_5_1; // @[RVTDNN.scala 72:63]
    outputReg_5_3 <= outputReg_5_2; // @[RVTDNN.scala 72:63]
    outputReg_5_4 <= outputReg_5_3; // @[RVTDNN.scala 72:63]
    outputReg_5_5 <= outputReg_5_4; // @[RVTDNN.scala 72:63]
    outputReg_6_0 <= BA_2_io_outAct_1; // @[RVTDNN.scala 73:63]
    outputReg_6_1 <= outputReg_6_0; // @[RVTDNN.scala 72:63]
    outputReg_6_2 <= outputReg_6_1; // @[RVTDNN.scala 72:63]
    outputReg_6_3 <= outputReg_6_2; // @[RVTDNN.scala 72:63]
    outputReg_6_4 <= outputReg_6_3; // @[RVTDNN.scala 72:63]
    outputReg_6_5 <= outputReg_6_4; // @[RVTDNN.scala 72:63]
    outputReg_6_6 <= outputReg_6_5; // @[RVTDNN.scala 72:63]
    outputReg_7_0 <= BA_2_io_outAct_0; // @[RVTDNN.scala 73:63]
    outputReg_7_1 <= outputReg_7_0; // @[RVTDNN.scala 72:63]
    outputReg_7_2 <= outputReg_7_1; // @[RVTDNN.scala 72:63]
    outputReg_7_3 <= outputReg_7_2; // @[RVTDNN.scala 72:63]
    outputReg_7_4 <= outputReg_7_3; // @[RVTDNN.scala 72:63]
    outputReg_7_5 <= outputReg_7_4; // @[RVTDNN.scala 72:63]
    outputReg_7_6 <= outputReg_7_5; // @[RVTDNN.scala 72:63]
    outputReg_7_7 <= outputReg_7_6; // @[RVTDNN.scala 72:63]
  end
endmodule
module RVTDNNTop(
  input         clock,
  input         reset,
  input  [15:0] io_bramIF_wrData,
  output [15:0] io_bramIF_rdData,
  input  [8:0]  io_bramIF_wrAddr,
  input  [8:0]  io_bramIF_rdAddr,
  input         io_bramIF_wrEn,
  input         io_load,
  input  [15:0] io_inAct_0,
  input  [15:0] io_inAct_1,
  input  [15:0] io_inAct_2,
  input  [15:0] io_inAct_3,
  input  [15:0] io_inAct_4,
  input  [15:0] io_inAct_5,
  input  [15:0] io_inAct_6,
  input  [15:0] io_inAct_7,
  output [15:0] io_outAct_0,
  output [15:0] io_outAct_1,
  output [15:0] io_outAct_2,
  output [15:0] io_outAct_3,
  output [15:0] io_outAct_4,
  output [15:0] io_outAct_5,
  output [15:0] io_outAct_6,
  output [15:0] io_outAct_7
);
  wire  loadModule_clock; // @[RVTDNNTop.scala 40:29]
  wire  loadModule_reset; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_bramIF_wrData; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_bramIF_rdData; // @[RVTDNNTop.scala 40:29]
  wire [8:0] loadModule_io_bramIF_wrAddr; // @[RVTDNNTop.scala 40:29]
  wire [8:0] loadModule_io_bramIF_rdAddr; // @[RVTDNNTop.scala 40:29]
  wire  loadModule_io_bramIF_wrEn; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_0; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_1; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_2; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_3; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_4; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_5; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_6; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_7; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_8; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outWeight_9; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_0; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_1; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_2; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_3; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_4; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_5; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_6; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_7; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_8; // @[RVTDNNTop.scala 40:29]
  wire [15:0] loadModule_io_outBias_9; // @[RVTDNNTop.scala 40:29]
  wire [2:0] loadModule_io_outWtValid; // @[RVTDNNTop.scala 40:29]
  wire [2:0] loadModule_io_outBiasValid; // @[RVTDNNTop.scala 40:29]
  wire  loadModule_io_load; // @[RVTDNNTop.scala 40:29]
  wire  rvtdnnModule_clock; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_0; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_1; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_2; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_3; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_4; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_5; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_6; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inAct_7; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_0; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_1; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_2; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_3; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_4; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_5; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_6; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_outAct_7; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_0; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_1; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_2; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_3; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_4; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_5; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_6; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_7; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_8; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inWeight_9; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_0; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_1; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_2; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_3; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_4; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_5; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_6; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_7; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_8; // @[RVTDNNTop.scala 42:29]
  wire [15:0] rvtdnnModule_io_inBias_9; // @[RVTDNNTop.scala 42:29]
  wire [2:0] rvtdnnModule_io_inWtValid; // @[RVTDNNTop.scala 42:29]
  wire [2:0] rvtdnnModule_io_inBiasValid; // @[RVTDNNTop.scala 42:29]
  LoadWeightBias loadModule ( // @[RVTDNNTop.scala 40:29]
    .clock(loadModule_clock),
    .reset(loadModule_reset),
    .io_bramIF_wrData(loadModule_io_bramIF_wrData),
    .io_bramIF_rdData(loadModule_io_bramIF_rdData),
    .io_bramIF_wrAddr(loadModule_io_bramIF_wrAddr),
    .io_bramIF_rdAddr(loadModule_io_bramIF_rdAddr),
    .io_bramIF_wrEn(loadModule_io_bramIF_wrEn),
    .io_outWeight_0(loadModule_io_outWeight_0),
    .io_outWeight_1(loadModule_io_outWeight_1),
    .io_outWeight_2(loadModule_io_outWeight_2),
    .io_outWeight_3(loadModule_io_outWeight_3),
    .io_outWeight_4(loadModule_io_outWeight_4),
    .io_outWeight_5(loadModule_io_outWeight_5),
    .io_outWeight_6(loadModule_io_outWeight_6),
    .io_outWeight_7(loadModule_io_outWeight_7),
    .io_outWeight_8(loadModule_io_outWeight_8),
    .io_outWeight_9(loadModule_io_outWeight_9),
    .io_outBias_0(loadModule_io_outBias_0),
    .io_outBias_1(loadModule_io_outBias_1),
    .io_outBias_2(loadModule_io_outBias_2),
    .io_outBias_3(loadModule_io_outBias_3),
    .io_outBias_4(loadModule_io_outBias_4),
    .io_outBias_5(loadModule_io_outBias_5),
    .io_outBias_6(loadModule_io_outBias_6),
    .io_outBias_7(loadModule_io_outBias_7),
    .io_outBias_8(loadModule_io_outBias_8),
    .io_outBias_9(loadModule_io_outBias_9),
    .io_outWtValid(loadModule_io_outWtValid),
    .io_outBiasValid(loadModule_io_outBiasValid),
    .io_load(loadModule_io_load)
  );
  RVTDNN rvtdnnModule ( // @[RVTDNNTop.scala 42:29]
    .clock(rvtdnnModule_clock),
    .io_inAct_0(rvtdnnModule_io_inAct_0),
    .io_inAct_1(rvtdnnModule_io_inAct_1),
    .io_inAct_2(rvtdnnModule_io_inAct_2),
    .io_inAct_3(rvtdnnModule_io_inAct_3),
    .io_inAct_4(rvtdnnModule_io_inAct_4),
    .io_inAct_5(rvtdnnModule_io_inAct_5),
    .io_inAct_6(rvtdnnModule_io_inAct_6),
    .io_inAct_7(rvtdnnModule_io_inAct_7),
    .io_outAct_0(rvtdnnModule_io_outAct_0),
    .io_outAct_1(rvtdnnModule_io_outAct_1),
    .io_outAct_2(rvtdnnModule_io_outAct_2),
    .io_outAct_3(rvtdnnModule_io_outAct_3),
    .io_outAct_4(rvtdnnModule_io_outAct_4),
    .io_outAct_5(rvtdnnModule_io_outAct_5),
    .io_outAct_6(rvtdnnModule_io_outAct_6),
    .io_outAct_7(rvtdnnModule_io_outAct_7),
    .io_inWeight_0(rvtdnnModule_io_inWeight_0),
    .io_inWeight_1(rvtdnnModule_io_inWeight_1),
    .io_inWeight_2(rvtdnnModule_io_inWeight_2),
    .io_inWeight_3(rvtdnnModule_io_inWeight_3),
    .io_inWeight_4(rvtdnnModule_io_inWeight_4),
    .io_inWeight_5(rvtdnnModule_io_inWeight_5),
    .io_inWeight_6(rvtdnnModule_io_inWeight_6),
    .io_inWeight_7(rvtdnnModule_io_inWeight_7),
    .io_inWeight_8(rvtdnnModule_io_inWeight_8),
    .io_inWeight_9(rvtdnnModule_io_inWeight_9),
    .io_inBias_0(rvtdnnModule_io_inBias_0),
    .io_inBias_1(rvtdnnModule_io_inBias_1),
    .io_inBias_2(rvtdnnModule_io_inBias_2),
    .io_inBias_3(rvtdnnModule_io_inBias_3),
    .io_inBias_4(rvtdnnModule_io_inBias_4),
    .io_inBias_5(rvtdnnModule_io_inBias_5),
    .io_inBias_6(rvtdnnModule_io_inBias_6),
    .io_inBias_7(rvtdnnModule_io_inBias_7),
    .io_inBias_8(rvtdnnModule_io_inBias_8),
    .io_inBias_9(rvtdnnModule_io_inBias_9),
    .io_inWtValid(rvtdnnModule_io_inWtValid),
    .io_inBiasValid(rvtdnnModule_io_inBiasValid)
  );
  assign io_bramIF_rdData = loadModule_io_bramIF_rdData; // @[RVTDNNTop.scala 56:29]
  assign io_outAct_0 = rvtdnnModule_io_outAct_0; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_1 = rvtdnnModule_io_outAct_1; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_2 = rvtdnnModule_io_outAct_2; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_3 = rvtdnnModule_io_outAct_3; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_4 = rvtdnnModule_io_outAct_4; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_5 = rvtdnnModule_io_outAct_5; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_6 = rvtdnnModule_io_outAct_6; // @[RVTDNNTop.scala 59:29]
  assign io_outAct_7 = rvtdnnModule_io_outAct_7; // @[RVTDNNTop.scala 59:29]
  assign loadModule_clock = clock;
  assign loadModule_reset = reset;
  assign loadModule_io_bramIF_wrData = io_bramIF_wrData; // @[RVTDNNTop.scala 56:29]
  assign loadModule_io_bramIF_wrAddr = io_bramIF_wrAddr; // @[RVTDNNTop.scala 56:29]
  assign loadModule_io_bramIF_rdAddr = io_bramIF_rdAddr; // @[RVTDNNTop.scala 56:29]
  assign loadModule_io_bramIF_wrEn = io_bramIF_wrEn; // @[RVTDNNTop.scala 56:29]
  assign loadModule_io_load = io_load; // @[RVTDNNTop.scala 57:29]
  assign rvtdnnModule_clock = clock;
  assign rvtdnnModule_io_inAct_0 = io_inAct_0; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_1 = io_inAct_1; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_2 = io_inAct_2; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_3 = io_inAct_3; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_4 = io_inAct_4; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_5 = io_inAct_5; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_6 = io_inAct_6; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inAct_7 = io_inAct_7; // @[RVTDNNTop.scala 58:29]
  assign rvtdnnModule_io_inWeight_0 = loadModule_io_outWeight_0; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_1 = loadModule_io_outWeight_1; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_2 = loadModule_io_outWeight_2; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_3 = loadModule_io_outWeight_3; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_4 = loadModule_io_outWeight_4; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_5 = loadModule_io_outWeight_5; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_6 = loadModule_io_outWeight_6; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_7 = loadModule_io_outWeight_7; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_8 = loadModule_io_outWeight_8; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inWeight_9 = loadModule_io_outWeight_9; // @[RVTDNNTop.scala 62:33]
  assign rvtdnnModule_io_inBias_0 = loadModule_io_outBias_0; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_1 = loadModule_io_outBias_1; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_2 = loadModule_io_outBias_2; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_3 = loadModule_io_outBias_3; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_4 = loadModule_io_outBias_4; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_5 = loadModule_io_outBias_5; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_6 = loadModule_io_outBias_6; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_7 = loadModule_io_outBias_7; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_8 = loadModule_io_outBias_8; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inBias_9 = loadModule_io_outBias_9; // @[RVTDNNTop.scala 63:33]
  assign rvtdnnModule_io_inWtValid = loadModule_io_outWtValid; // @[RVTDNNTop.scala 64:33]
  assign rvtdnnModule_io_inBiasValid = loadModule_io_outBiasValid; // @[RVTDNNTop.scala 65:33]
endmodule
